
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity start_menu is
--FPGA pin decleration
    Port (	clk			:  in std_logic;
				reset			:  in std_logic;
				x_counter   :  in integer range 0 to 640;
				y_counter	:	in integer range 0 to 480;
				RGB    		: 	out STD_LOGIC_VECTOR(2 downto 0));  --VGA RGB output
				
end start_menu;

architecture Behavioral of start_menu is

    signal animation_on : std_logic; --flashing the "PRESS ANY KEY"
begin

-------------------------------------------Animation-----------------------------------------------------
    process(clk,reset)
        variable    animation_timer_var : integer range 0 to 25000000;
        begin
            if(reset = '1') then
                animation_timer_var := 0;
                animation_on <= '0';
                
            elsif (clk'event and clk = '1') then
                animation_timer_var := animation_timer_var + 1;
                    if(animation_timer_var = 25000000) then
                        animation_timer_var := 0;
                        animation_on <= not(animation_on);
                    end if;
            end if;
        
        end process;

    RGB			  <= "111" when  		( y_counter = 98 AND ((x_counter >= 172 AND x_counter <= 197 ) ))
											OR ( y_counter = 99 AND ((x_counter >= 172 AND x_counter <= 197 ) ))
											OR ( y_counter = 100 AND ((x_counter >= 172 AND x_counter <= 197 ) ))
											OR ( y_counter = 101 AND ((x_counter >= 172 AND x_counter <= 197 ) ))
											OR ( y_counter = 102 AND ((x_counter >= 172 AND x_counter <= 197 ) ))
											OR ( y_counter = 103 AND ((x_counter >= 172 AND x_counter <= 197 ) ))
											OR ( y_counter = 104 AND ((x_counter >= 172 AND x_counter <= 197 ) OR (x_counter >= 344 AND x_counter <= 360 ) ))
											OR ( y_counter = 105 AND ((x_counter >= 172 AND x_counter <= 197 ) OR (x_counter >= 344 AND x_counter <= 360 ) ))
											OR ( y_counter = 106 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 192 AND x_counter <= 202 ) OR (x_counter >= 344 AND x_counter <= 360 ) ))
											OR ( y_counter = 107 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 192 AND x_counter <= 202 ) OR (x_counter >= 344 AND x_counter <= 360 ) ))
											OR ( y_counter = 108 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 192 AND x_counter <= 202 ) OR (x_counter >= 340 AND x_counter <= 348 ) OR (x_counter >= 356 AND x_counter <= 364 ) ))
											OR ( y_counter = 109 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 192 AND x_counter <= 202 ) OR (x_counter >= 340 AND x_counter <= 348 ) OR (x_counter >= 356 AND x_counter <= 364 ) ))
											OR ( y_counter = 110 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 192 AND x_counter <= 202 ) OR (x_counter >= 340 AND x_counter <= 348 ) OR (x_counter >= 356 AND x_counter <= 364 ) ))
											OR ( y_counter = 111 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 192 AND x_counter <= 202 ) OR (x_counter >= 340 AND x_counter <= 348 ) OR (x_counter >= 356 AND x_counter <= 364 ) ))
											OR ( y_counter = 112 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 192 AND x_counter <= 202 ) OR (x_counter >= 216 AND x_counter <= 232 ) OR (x_counter >= 244 AND x_counter <= 264 ) OR (x_counter >= 280 AND x_counter <= 300 ) OR (x_counter >= 340 AND x_counter <= 348 ) OR (x_counter >= 356 AND x_counter <= 364 ) OR (x_counter >= 376 AND x_counter <= 392 ) OR (x_counter >= 404 AND x_counter <= 428 ) OR (x_counter >= 440 AND x_counter <= 456 ) ))
											OR ( y_counter = 113 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 192 AND x_counter <= 202 ) OR (x_counter >= 216 AND x_counter <= 232 ) OR (x_counter >= 244 AND x_counter <= 264 ) OR (x_counter >= 280 AND x_counter <= 300 ) OR (x_counter >= 340 AND x_counter <= 348 ) OR (x_counter >= 356 AND x_counter <= 364 ) OR (x_counter >= 376 AND x_counter <= 392 ) OR (x_counter >= 404 AND x_counter <= 428 ) OR (x_counter >= 440 AND x_counter <= 456 ) ))
											OR ( y_counter = 114 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 192 AND x_counter <= 202 ) OR (x_counter >= 216 AND x_counter <= 232 ) OR (x_counter >= 244 AND x_counter <= 264 ) OR (x_counter >= 280 AND x_counter <= 300 ) OR (x_counter >= 340 AND x_counter <= 348 ) OR (x_counter >= 356 AND x_counter <= 364 ) OR (x_counter >= 376 AND x_counter <= 392 ) OR (x_counter >= 404 AND x_counter <= 428 ) OR (x_counter >= 440 AND x_counter <= 456 ) ))
											OR ( y_counter = 115 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 192 AND x_counter <= 202 ) OR (x_counter >= 216 AND x_counter <= 232 ) OR (x_counter >= 244 AND x_counter <= 264 ) OR (x_counter >= 280 AND x_counter <= 300 ) OR (x_counter >= 340 AND x_counter <= 348 ) OR (x_counter >= 356 AND x_counter <= 364 ) OR (x_counter >= 376 AND x_counter <= 392 ) OR (x_counter >= 404 AND x_counter <= 428 ) OR (x_counter >= 440 AND x_counter <= 456 ) ))
											OR ( y_counter = 116 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 192 AND x_counter <= 202 ) OR (x_counter >= 212 AND x_counter <= 220 ) OR (x_counter >= 228 AND x_counter <= 236 ) OR (x_counter >= 244 AND x_counter <= 252 ) OR (x_counter >= 260 AND x_counter <= 268 ) OR (x_counter >= 276 AND x_counter <= 284 ) OR (x_counter >= 292 AND x_counter <= 300 ) OR (x_counter >= 340 AND x_counter <= 348 ) OR (x_counter >= 388 AND x_counter <= 396 ) OR (x_counter >= 404 AND x_counter <= 412 ) OR (x_counter >= 416 AND x_counter <= 420 ) OR (x_counter >= 424 AND x_counter <= 432 ) OR (x_counter >= 436 AND x_counter <= 444 ) OR (x_counter >= 452 AND x_counter <= 460 ) ))
											OR ( y_counter = 117 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 192 AND x_counter <= 202 ) OR (x_counter >= 212 AND x_counter <= 220 ) OR (x_counter >= 228 AND x_counter <= 236 ) OR (x_counter >= 244 AND x_counter <= 252 ) OR (x_counter >= 260 AND x_counter <= 268 ) OR (x_counter >= 276 AND x_counter <= 284 ) OR (x_counter >= 292 AND x_counter <= 300 ) OR (x_counter >= 340 AND x_counter <= 348 ) OR (x_counter >= 388 AND x_counter <= 396 ) OR (x_counter >= 404 AND x_counter <= 412 ) OR (x_counter >= 416 AND x_counter <= 420 ) OR (x_counter >= 424 AND x_counter <= 432 ) OR (x_counter >= 436 AND x_counter <= 444 ) OR (x_counter >= 452 AND x_counter <= 460 ) ))
											OR ( y_counter = 118 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 192 AND x_counter <= 202 ) OR (x_counter >= 212 AND x_counter <= 220 ) OR (x_counter >= 228 AND x_counter <= 236 ) OR (x_counter >= 244 AND x_counter <= 252 ) OR (x_counter >= 260 AND x_counter <= 268 ) OR (x_counter >= 276 AND x_counter <= 284 ) OR (x_counter >= 292 AND x_counter <= 300 ) OR (x_counter >= 340 AND x_counter <= 348 ) OR (x_counter >= 388 AND x_counter <= 396 ) OR (x_counter >= 404 AND x_counter <= 412 ) OR (x_counter >= 416 AND x_counter <= 420 ) OR (x_counter >= 424 AND x_counter <= 432 ) OR (x_counter >= 436 AND x_counter <= 444 ) OR (x_counter >= 452 AND x_counter <= 460 ) ))
											OR ( y_counter = 119 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 192 AND x_counter <= 202 ) OR (x_counter >= 212 AND x_counter <= 220 ) OR (x_counter >= 228 AND x_counter <= 236 ) OR (x_counter >= 244 AND x_counter <= 252 ) OR (x_counter >= 260 AND x_counter <= 268 ) OR (x_counter >= 276 AND x_counter <= 284 ) OR (x_counter >= 292 AND x_counter <= 300 ) OR (x_counter >= 340 AND x_counter <= 348 ) OR (x_counter >= 388 AND x_counter <= 396 ) OR (x_counter >= 404 AND x_counter <= 412 ) OR (x_counter >= 416 AND x_counter <= 420 ) OR (x_counter >= 424 AND x_counter <= 432 ) OR (x_counter >= 436 AND x_counter <= 444 ) OR (x_counter >= 452 AND x_counter <= 460 ) ))
											OR ( y_counter = 120 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 192 AND x_counter <= 202 ) OR (x_counter >= 212 AND x_counter <= 220 ) OR (x_counter >= 228 AND x_counter <= 236 ) OR (x_counter >= 244 AND x_counter <= 252 ) OR (x_counter >= 260 AND x_counter <= 268 ) OR (x_counter >= 276 AND x_counter <= 284 ) OR (x_counter >= 292 AND x_counter <= 300 ) OR (x_counter >= 340 AND x_counter <= 348 ) OR (x_counter >= 388 AND x_counter <= 396 ) OR (x_counter >= 404 AND x_counter <= 412 ) OR (x_counter >= 416 AND x_counter <= 420 ) OR (x_counter >= 424 AND x_counter <= 432 ) OR (x_counter >= 436 AND x_counter <= 444 ) OR (x_counter >= 452 AND x_counter <= 460 ) ))
											OR ( y_counter = 121 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 192 AND x_counter <= 202 ) OR (x_counter >= 212 AND x_counter <= 220 ) OR (x_counter >= 228 AND x_counter <= 236 ) OR (x_counter >= 244 AND x_counter <= 252 ) OR (x_counter >= 260 AND x_counter <= 268 ) OR (x_counter >= 276 AND x_counter <= 284 ) OR (x_counter >= 292 AND x_counter <= 300 ) OR (x_counter >= 340 AND x_counter <= 348 ) OR (x_counter >= 388 AND x_counter <= 396 ) OR (x_counter >= 404 AND x_counter <= 412 ) OR (x_counter >= 416 AND x_counter <= 420 ) OR (x_counter >= 424 AND x_counter <= 432 ) OR (x_counter >= 436 AND x_counter <= 444 ) OR (x_counter >= 452 AND x_counter <= 460 ) ))
											OR ( y_counter = 122 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 192 AND x_counter <= 202 ) OR (x_counter >= 212 AND x_counter <= 220 ) OR (x_counter >= 228 AND x_counter <= 236 ) OR (x_counter >= 244 AND x_counter <= 252 ) OR (x_counter >= 260 AND x_counter <= 268 ) OR (x_counter >= 276 AND x_counter <= 284 ) OR (x_counter >= 292 AND x_counter <= 300 ) OR (x_counter >= 340 AND x_counter <= 348 ) OR (x_counter >= 388 AND x_counter <= 396 ) OR (x_counter >= 404 AND x_counter <= 412 ) OR (x_counter >= 416 AND x_counter <= 420 ) OR (x_counter >= 424 AND x_counter <= 432 ) OR (x_counter >= 436 AND x_counter <= 444 ) OR (x_counter >= 452 AND x_counter <= 460 ) ))
											OR ( y_counter = 123 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 192 AND x_counter <= 202 ) OR (x_counter >= 212 AND x_counter <= 220 ) OR (x_counter >= 228 AND x_counter <= 236 ) OR (x_counter >= 244 AND x_counter <= 252 ) OR (x_counter >= 260 AND x_counter <= 268 ) OR (x_counter >= 276 AND x_counter <= 284 ) OR (x_counter >= 292 AND x_counter <= 300 ) OR (x_counter >= 340 AND x_counter <= 348 ) OR (x_counter >= 388 AND x_counter <= 396 ) OR (x_counter >= 404 AND x_counter <= 412 ) OR (x_counter >= 416 AND x_counter <= 420 ) OR (x_counter >= 424 AND x_counter <= 432 ) OR (x_counter >= 436 AND x_counter <= 444 ) OR (x_counter >= 452 AND x_counter <= 460 ) ))
											OR ( y_counter = 124 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 192 AND x_counter <= 202 ) OR (x_counter >= 212 AND x_counter <= 220 ) OR (x_counter >= 228 AND x_counter <= 236 ) OR (x_counter >= 244 AND x_counter <= 252 ) OR (x_counter >= 260 AND x_counter <= 268 ) OR (x_counter >= 276 AND x_counter <= 284 ) OR (x_counter >= 292 AND x_counter <= 300 ) OR (x_counter >= 340 AND x_counter <= 348 ) OR (x_counter >= 352 AND x_counter <= 364 ) OR (x_counter >= 376 AND x_counter <= 396 ) OR (x_counter >= 404 AND x_counter <= 412 ) OR (x_counter >= 416 AND x_counter <= 420 ) OR (x_counter >= 424 AND x_counter <= 432 ) OR (x_counter >= 436 AND x_counter <= 460 ) ))
											OR ( y_counter = 125 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 192 AND x_counter <= 202 ) OR (x_counter >= 212 AND x_counter <= 220 ) OR (x_counter >= 228 AND x_counter <= 236 ) OR (x_counter >= 244 AND x_counter <= 252 ) OR (x_counter >= 260 AND x_counter <= 268 ) OR (x_counter >= 276 AND x_counter <= 284 ) OR (x_counter >= 292 AND x_counter <= 300 ) OR (x_counter >= 340 AND x_counter <= 348 ) OR (x_counter >= 352 AND x_counter <= 364 ) OR (x_counter >= 376 AND x_counter <= 396 ) OR (x_counter >= 404 AND x_counter <= 412 ) OR (x_counter >= 416 AND x_counter <= 420 ) OR (x_counter >= 424 AND x_counter <= 432 ) OR (x_counter >= 436 AND x_counter <= 460 ) ))
											OR ( y_counter = 126 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 192 AND x_counter <= 202 ) OR (x_counter >= 212 AND x_counter <= 220 ) OR (x_counter >= 228 AND x_counter <= 236 ) OR (x_counter >= 244 AND x_counter <= 252 ) OR (x_counter >= 260 AND x_counter <= 268 ) OR (x_counter >= 276 AND x_counter <= 284 ) OR (x_counter >= 292 AND x_counter <= 300 ) OR (x_counter >= 340 AND x_counter <= 348 ) OR (x_counter >= 352 AND x_counter <= 364 ) OR (x_counter >= 376 AND x_counter <= 396 ) OR (x_counter >= 404 AND x_counter <= 412 ) OR (x_counter >= 416 AND x_counter <= 420 ) OR (x_counter >= 424 AND x_counter <= 432 ) OR (x_counter >= 436 AND x_counter <= 460 ) ))
											OR ( y_counter = 127 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 192 AND x_counter <= 202 ) OR (x_counter >= 212 AND x_counter <= 220 ) OR (x_counter >= 228 AND x_counter <= 236 ) OR (x_counter >= 244 AND x_counter <= 252 ) OR (x_counter >= 260 AND x_counter <= 268 ) OR (x_counter >= 276 AND x_counter <= 284 ) OR (x_counter >= 292 AND x_counter <= 300 ) OR (x_counter >= 340 AND x_counter <= 348 ) OR (x_counter >= 352 AND x_counter <= 364 ) OR (x_counter >= 376 AND x_counter <= 396 ) OR (x_counter >= 404 AND x_counter <= 412 ) OR (x_counter >= 416 AND x_counter <= 420 ) OR (x_counter >= 424 AND x_counter <= 432 ) OR (x_counter >= 436 AND x_counter <= 460 ) ))
											OR ( y_counter = 128 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 192 AND x_counter <= 202 ) OR (x_counter >= 212 AND x_counter <= 220 ) OR (x_counter >= 228 AND x_counter <= 236 ) OR (x_counter >= 244 AND x_counter <= 252 ) OR (x_counter >= 260 AND x_counter <= 268 ) OR (x_counter >= 276 AND x_counter <= 284 ) OR (x_counter >= 292 AND x_counter <= 300 ) OR (x_counter >= 340 AND x_counter <= 348 ) OR (x_counter >= 356 AND x_counter <= 364 ) OR (x_counter >= 372 AND x_counter <= 380 ) OR (x_counter >= 388 AND x_counter <= 396 ) OR (x_counter >= 404 AND x_counter <= 412 ) OR (x_counter >= 416 AND x_counter <= 420 ) OR (x_counter >= 424 AND x_counter <= 432 ) OR (x_counter >= 436 AND x_counter <= 444 ) ))
											OR ( y_counter = 129 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 192 AND x_counter <= 202 ) OR (x_counter >= 212 AND x_counter <= 220 ) OR (x_counter >= 228 AND x_counter <= 236 ) OR (x_counter >= 244 AND x_counter <= 252 ) OR (x_counter >= 260 AND x_counter <= 268 ) OR (x_counter >= 276 AND x_counter <= 284 ) OR (x_counter >= 292 AND x_counter <= 300 ) OR (x_counter >= 340 AND x_counter <= 348 ) OR (x_counter >= 356 AND x_counter <= 364 ) OR (x_counter >= 372 AND x_counter <= 380 ) OR (x_counter >= 388 AND x_counter <= 396 ) OR (x_counter >= 404 AND x_counter <= 412 ) OR (x_counter >= 416 AND x_counter <= 420 ) OR (x_counter >= 424 AND x_counter <= 432 ) OR (x_counter >= 436 AND x_counter <= 444 ) ))
											OR ( y_counter = 130 AND ((x_counter >= 172 AND x_counter <= 197 ) OR (x_counter >= 212 AND x_counter <= 220 ) OR (x_counter >= 228 AND x_counter <= 236 ) OR (x_counter >= 244 AND x_counter <= 252 ) OR (x_counter >= 260 AND x_counter <= 268 ) OR (x_counter >= 276 AND x_counter <= 284 ) OR (x_counter >= 292 AND x_counter <= 300 ) OR (x_counter >= 340 AND x_counter <= 348 ) OR (x_counter >= 356 AND x_counter <= 364 ) OR (x_counter >= 372 AND x_counter <= 380 ) OR (x_counter >= 388 AND x_counter <= 396 ) OR (x_counter >= 404 AND x_counter <= 412 ) OR (x_counter >= 416 AND x_counter <= 420 ) OR (x_counter >= 424 AND x_counter <= 432 ) OR (x_counter >= 436 AND x_counter <= 444 ) ))
											OR ( y_counter = 131 AND ((x_counter >= 172 AND x_counter <= 197 ) OR (x_counter >= 212 AND x_counter <= 220 ) OR (x_counter >= 228 AND x_counter <= 236 ) OR (x_counter >= 244 AND x_counter <= 252 ) OR (x_counter >= 260 AND x_counter <= 268 ) OR (x_counter >= 276 AND x_counter <= 284 ) OR (x_counter >= 292 AND x_counter <= 300 ) OR (x_counter >= 340 AND x_counter <= 348 ) OR (x_counter >= 356 AND x_counter <= 364 ) OR (x_counter >= 372 AND x_counter <= 380 ) OR (x_counter >= 388 AND x_counter <= 396 ) OR (x_counter >= 404 AND x_counter <= 412 ) OR (x_counter >= 416 AND x_counter <= 420 ) OR (x_counter >= 424 AND x_counter <= 432 ) OR (x_counter >= 436 AND x_counter <= 444 ) ))
											OR ( y_counter = 132 AND ((x_counter >= 172 AND x_counter <= 197 ) OR (x_counter >= 212 AND x_counter <= 220 ) OR (x_counter >= 228 AND x_counter <= 236 ) OR (x_counter >= 244 AND x_counter <= 252 ) OR (x_counter >= 260 AND x_counter <= 268 ) OR (x_counter >= 276 AND x_counter <= 284 ) OR (x_counter >= 292 AND x_counter <= 300 ) OR (x_counter >= 340 AND x_counter <= 348 ) OR (x_counter >= 356 AND x_counter <= 364 ) OR (x_counter >= 372 AND x_counter <= 380 ) OR (x_counter >= 388 AND x_counter <= 396 ) OR (x_counter >= 404 AND x_counter <= 412 ) OR (x_counter >= 416 AND x_counter <= 420 ) OR (x_counter >= 424 AND x_counter <= 432 ) OR (x_counter >= 436 AND x_counter <= 444 ) ))
											OR ( y_counter = 133 AND ((x_counter >= 172 AND x_counter <= 197 ) OR (x_counter >= 212 AND x_counter <= 220 ) OR (x_counter >= 228 AND x_counter <= 236 ) OR (x_counter >= 244 AND x_counter <= 252 ) OR (x_counter >= 260 AND x_counter <= 268 ) OR (x_counter >= 276 AND x_counter <= 284 ) OR (x_counter >= 292 AND x_counter <= 300 ) OR (x_counter >= 340 AND x_counter <= 348 ) OR (x_counter >= 356 AND x_counter <= 364 ) OR (x_counter >= 372 AND x_counter <= 380 ) OR (x_counter >= 388 AND x_counter <= 396 ) OR (x_counter >= 404 AND x_counter <= 412 ) OR (x_counter >= 416 AND x_counter <= 420 ) OR (x_counter >= 424 AND x_counter <= 432 ) OR (x_counter >= 436 AND x_counter <= 444 ) ))
											OR ( y_counter = 134 AND ((x_counter >= 172 AND x_counter <= 197 ) OR (x_counter >= 212 AND x_counter <= 220 ) OR (x_counter >= 228 AND x_counter <= 236 ) OR (x_counter >= 244 AND x_counter <= 252 ) OR (x_counter >= 260 AND x_counter <= 268 ) OR (x_counter >= 276 AND x_counter <= 284 ) OR (x_counter >= 292 AND x_counter <= 300 ) OR (x_counter >= 340 AND x_counter <= 348 ) OR (x_counter >= 356 AND x_counter <= 364 ) OR (x_counter >= 372 AND x_counter <= 380 ) OR (x_counter >= 388 AND x_counter <= 396 ) OR (x_counter >= 404 AND x_counter <= 412 ) OR (x_counter >= 416 AND x_counter <= 420 ) OR (x_counter >= 424 AND x_counter <= 432 ) OR (x_counter >= 436 AND x_counter <= 444 ) ))
											OR ( y_counter = 135 AND ((x_counter >= 172 AND x_counter <= 197 ) OR (x_counter >= 212 AND x_counter <= 220 ) OR (x_counter >= 228 AND x_counter <= 236 ) OR (x_counter >= 244 AND x_counter <= 252 ) OR (x_counter >= 260 AND x_counter <= 268 ) OR (x_counter >= 276 AND x_counter <= 284 ) OR (x_counter >= 292 AND x_counter <= 300 ) OR (x_counter >= 340 AND x_counter <= 348 ) OR (x_counter >= 356 AND x_counter <= 364 ) OR (x_counter >= 372 AND x_counter <= 380 ) OR (x_counter >= 388 AND x_counter <= 396 ) OR (x_counter >= 404 AND x_counter <= 412 ) OR (x_counter >= 416 AND x_counter <= 420 ) OR (x_counter >= 424 AND x_counter <= 432 ) OR (x_counter >= 436 AND x_counter <= 444 ) ))
											OR ( y_counter = 136 AND ((x_counter >= 172 AND x_counter <= 197 ) OR (x_counter >= 216 AND x_counter <= 232 ) OR (x_counter >= 244 AND x_counter <= 252 ) OR (x_counter >= 260 AND x_counter <= 268 ) OR (x_counter >= 280 AND x_counter <= 300 ) OR (x_counter >= 344 AND x_counter <= 364 ) OR (x_counter >= 376 AND x_counter <= 396 ) OR (x_counter >= 404 AND x_counter <= 412 ) OR (x_counter >= 424 AND x_counter <= 432 ) OR (x_counter >= 440 AND x_counter <= 456 ) ))
											OR ( y_counter = 137 AND ((x_counter >= 172 AND x_counter <= 197 ) OR (x_counter >= 216 AND x_counter <= 232 ) OR (x_counter >= 244 AND x_counter <= 252 ) OR (x_counter >= 260 AND x_counter <= 268 ) OR (x_counter >= 280 AND x_counter <= 300 ) OR (x_counter >= 344 AND x_counter <= 364 ) OR (x_counter >= 376 AND x_counter <= 396 ) OR (x_counter >= 404 AND x_counter <= 412 ) OR (x_counter >= 424 AND x_counter <= 432 ) OR (x_counter >= 440 AND x_counter <= 456 ) ))
											OR ( y_counter = 138 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 216 AND x_counter <= 232 ) OR (x_counter >= 244 AND x_counter <= 252 ) OR (x_counter >= 260 AND x_counter <= 268 ) OR (x_counter >= 280 AND x_counter <= 300 ) OR (x_counter >= 344 AND x_counter <= 364 ) OR (x_counter >= 376 AND x_counter <= 396 ) OR (x_counter >= 404 AND x_counter <= 412 ) OR (x_counter >= 424 AND x_counter <= 432 ) OR (x_counter >= 440 AND x_counter <= 456 ) ))
											OR ( y_counter = 139 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 216 AND x_counter <= 232 ) OR (x_counter >= 244 AND x_counter <= 252 ) OR (x_counter >= 260 AND x_counter <= 268 ) OR (x_counter >= 280 AND x_counter <= 300 ) OR (x_counter >= 344 AND x_counter <= 364 ) OR (x_counter >= 376 AND x_counter <= 396 ) OR (x_counter >= 404 AND x_counter <= 412 ) OR (x_counter >= 424 AND x_counter <= 432 ) OR (x_counter >= 440 AND x_counter <= 456 ) ))
											OR ( y_counter = 140 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 292 AND x_counter <= 300 ) ))
											OR ( y_counter = 141 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 292 AND x_counter <= 300 ) ))
											OR ( y_counter = 142 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 292 AND x_counter <= 300 ) ))
											OR ( y_counter = 143 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 292 AND x_counter <= 300 ) ))
											OR ( y_counter = 144 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 292 AND x_counter <= 300 ) ))
											OR ( y_counter = 145 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 292 AND x_counter <= 300 ) ))
											OR ( y_counter = 146 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 292 AND x_counter <= 300 ) ))
											OR ( y_counter = 147 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 292 AND x_counter <= 300 ) ))
											OR ( y_counter = 148 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 276 AND x_counter <= 296 ) ))
											OR ( y_counter = 149 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 276 AND x_counter <= 296 ) ))
											OR ( y_counter = 150 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 276 AND x_counter <= 296 ) ))
											OR ( y_counter = 151 AND ((x_counter >= 172 AND x_counter <= 182 ) OR (x_counter >= 276 AND x_counter <= 296 ) ))
											OR ( y_counter = 152 AND ((x_counter >= 172 AND x_counter <= 182 ) ))
											OR ( y_counter = 153 AND ((x_counter >= 172 AND x_counter <= 182 ) ))
											OR ( y_counter = 154 AND ((x_counter >= 172 AND x_counter <= 182 ) ))
											OR ( y_counter = 155 AND ((x_counter >= 172 AND x_counter <= 182 ) ))
											OR ( y_counter = 156 AND ((x_counter >= 172 AND x_counter <= 182 ) ))
											OR ( y_counter = 157 AND ((x_counter >= 172 AND x_counter <= 182 ) ))
											OR ( y_counter = 158 AND ((x_counter >= 172 AND x_counter <= 182 ) ))
											OR ( y_counter = 159 AND ((x_counter >= 172 AND x_counter <= 182 ) ))
											OR ( y_counter = 160 AND ((x_counter >= 172 AND x_counter <= 182 ) ))
											OR ( y_counter = 161 AND ((x_counter >= 172 AND x_counter <= 182 ) ))
											OR ( y_counter = 162 AND ((x_counter >= 172 AND x_counter <= 182 ) ))
											OR ( y_counter = 163 AND ((x_counter >= 172 AND x_counter <= 182 ) ))
											OR ( y_counter = 164 AND ((x_counter >= 172 AND x_counter <= 182 ) ))
											OR ( y_counter = 165 AND ((x_counter >= 172 AND x_counter <= 182 ) ))
											OR ( y_counter = 166 AND ((x_counter >= 172 AND x_counter <= 182 ) ))
											OR ( y_counter = 167 AND ((x_counter >= 172 AND x_counter <= 182 ) ))
											OR ( y_counter = 168 AND ((x_counter >= 172 AND x_counter <= 182 ) ))
											OR ( y_counter = 169 AND ((x_counter >= 172 AND x_counter <= 182 ) ))
											OR ( y_counter = 220 AND animation_on ='1' AND ((x_counter >= 267 AND x_counter <= 272 ) OR (x_counter >= 316 AND x_counter <= 320 ) OR (x_counter >= 324 AND x_counter <= 326 ) OR (x_counter >= 348 AND x_counter <= 350 ) )) --START ANIMATION
											OR ( y_counter = 221 AND animation_on ='1' AND ((x_counter >= 267 AND x_counter <= 269 ) OR (x_counter >= 271 AND x_counter <= 273 ) OR (x_counter >= 315 AND x_counter <= 317 ) OR (x_counter >= 319 AND x_counter <= 321 ) OR (x_counter >= 324 AND x_counter <= 326 ) OR (x_counter >= 348 AND x_counter <= 350 ) ))
											OR ( y_counter = 222 AND animation_on ='1' AND ((x_counter >= 267 AND x_counter <= 269 ) OR (x_counter >= 271 AND x_counter <= 273 ) OR (x_counter >= 275 AND x_counter <= 277 ) OR (x_counter >= 279 AND x_counter <= 281 ) OR (x_counter >= 284 AND x_counter <= 288 ) OR (x_counter >= 292 AND x_counter <= 297 ) OR (x_counter >= 300 AND x_counter <= 305 ) OR (x_counter >= 315 AND x_counter <= 317 ) OR (x_counter >= 323 AND x_counter <= 329 ) OR (x_counter >= 332 AND x_counter <= 336 ) OR (x_counter >= 339 AND x_counter <= 341 ) OR (x_counter >= 343 AND x_counter <= 345 ) OR (x_counter >= 347 AND x_counter <= 353 ) ))
											OR ( y_counter = 223 AND animation_on ='1' AND ((x_counter >= 267 AND x_counter <= 269 ) OR (x_counter >= 271 AND x_counter <= 273 ) OR (x_counter >= 275 AND x_counter <= 277 ) OR (x_counter >= 278 AND x_counter <= 281 ) OR (x_counter >= 283 AND x_counter <= 285 ) OR (x_counter >= 287 AND x_counter <= 289 ) OR (x_counter >= 291 AND x_counter <= 293 ) OR (x_counter >= 299 AND x_counter <= 301 ) OR (x_counter >= 316 AND x_counter <= 318 ) OR (x_counter >= 324 AND x_counter <= 326 ) OR (x_counter >= 335 AND x_counter <= 337 ) OR (x_counter >= 339 AND x_counter <= 341 ) OR (x_counter >= 342 AND x_counter <= 345 ) OR (x_counter >= 348 AND x_counter <= 350 ) ))
											OR ( y_counter = 224 AND animation_on ='1' AND ((x_counter >= 267 AND x_counter <= 272 ) OR (x_counter >= 275 AND x_counter <= 278 ) OR (x_counter >= 283 AND x_counter <= 285 ) OR (x_counter >= 287 AND x_counter <= 289 ) OR (x_counter >= 291 AND x_counter <= 293 ) OR (x_counter >= 299 AND x_counter <= 301 ) OR (x_counter >= 317 AND x_counter <= 319 ) OR (x_counter >= 324 AND x_counter <= 326 ) OR (x_counter >= 335 AND x_counter <= 337 ) OR (x_counter >= 339 AND x_counter <= 342 ) OR (x_counter >= 348 AND x_counter <= 350 ) ))
											OR ( y_counter = 225 AND animation_on ='1' AND ((x_counter >= 267 AND x_counter <= 269 ) OR (x_counter >= 275 AND x_counter <= 277 ) OR (x_counter >= 283 AND x_counter <= 289 ) OR (x_counter >= 292 AND x_counter <= 296 ) OR (x_counter >= 300 AND x_counter <= 304 ) OR (x_counter >= 318 AND x_counter <= 320 ) OR (x_counter >= 324 AND x_counter <= 326 ) OR (x_counter >= 332 AND x_counter <= 337 ) OR (x_counter >= 339 AND x_counter <= 341 ) OR (x_counter >= 348 AND x_counter <= 350 ) ))
											OR ( y_counter = 226 AND animation_on ='1' AND ((x_counter >= 267 AND x_counter <= 269 ) OR (x_counter >= 275 AND x_counter <= 277 ) OR (x_counter >= 283 AND x_counter <= 285 ) OR (x_counter >= 295 AND x_counter <= 297 ) OR (x_counter >= 303 AND x_counter <= 305 ) OR (x_counter >= 319 AND x_counter <= 321 ) OR (x_counter >= 324 AND x_counter <= 326 ) OR (x_counter >= 331 AND x_counter <= 333 ) OR (x_counter >= 335 AND x_counter <= 337 ) OR (x_counter >= 339 AND x_counter <= 341 ) OR (x_counter >= 348 AND x_counter <= 350 ) ))
											OR ( y_counter = 227 AND animation_on ='1' AND ((x_counter >= 267 AND x_counter <= 269 ) OR (x_counter >= 275 AND x_counter <= 277 ) OR (x_counter >= 283 AND x_counter <= 285 ) OR (x_counter >= 295 AND x_counter <= 297 ) OR (x_counter >= 303 AND x_counter <= 305 ) OR (x_counter >= 315 AND x_counter <= 317 ) OR (x_counter >= 319 AND x_counter <= 321 ) OR (x_counter >= 324 AND x_counter <= 326 ) OR (x_counter >= 331 AND x_counter <= 333 ) OR (x_counter >= 335 AND x_counter <= 337 ) OR (x_counter >= 339 AND x_counter <= 341 ) OR (x_counter >= 348 AND x_counter <= 350 ) ))
											OR ( y_counter = 228 AND animation_on ='1' AND ((x_counter >= 267 AND x_counter <= 269 ) OR (x_counter >= 275 AND x_counter <= 277 ) OR (x_counter >= 284 AND x_counter <= 288 ) OR (x_counter >= 291 AND x_counter <= 296 ) OR (x_counter >= 299 AND x_counter <= 304 ) OR (x_counter >= 316 AND x_counter <= 320 ) OR (x_counter >= 325 AND x_counter <= 329 ) OR (x_counter >= 332 AND x_counter <= 337 ) OR (x_counter >= 339 AND x_counter <= 341 ) OR (x_counter >= 349 AND x_counter <= 353 ) )) --END ANIMATION


											OR	(y_counter = 362 AND ((x_counter >= 208 AND x_counter <= 225) OR (x_counter >= 229 AND x_counter <= 234) OR (x_counter >= 238 AND x_counter <= 243) OR (x_counter >= 325 AND x_counter <= 342) OR (x_counter >= 346 AND x_counter <= 351) OR (x_counter >= 355 AND x_counter <= 360) OR (x_counter >= 848 AND x_counter <= 865) OR (x_counter >= 869 AND x_counter <= 874) OR (x_counter >= 878 AND x_counter <= 883) OR (x_counter >= 965 AND x_counter <= 982) OR (x_counter >= 986 AND x_counter <= 991) OR (x_counter >= 995 AND x_counter <= 1000) OR (x_counter >= 1488 AND x_counter <= 1505) OR (x_counter >= 1509 AND x_counter <= 1514) OR (x_counter >= 1518 AND x_counter <= 1523) OR (x_counter >= 1605 AND x_counter <= 1622) OR (x_counter >= 1626 AND x_counter <= 1631) OR (x_counter >= 1635 AND x_counter <= 1640)))
											OR	(y_counter = 363 AND ((x_counter >= 208 AND x_counter <= 225) OR (x_counter >= 229 AND x_counter <= 234) OR (x_counter >= 238 AND x_counter <= 243) OR (x_counter >= 325 AND x_counter <= 342) OR (x_counter >= 346 AND x_counter <= 351) OR (x_counter >= 355 AND x_counter <= 360) OR (x_counter >= 848 AND x_counter <= 865) OR (x_counter >= 869 AND x_counter <= 874) OR (x_counter >= 878 AND x_counter <= 883) OR (x_counter >= 965 AND x_counter <= 982) OR (x_counter >= 986 AND x_counter <= 991) OR (x_counter >= 995 AND x_counter <= 1000) OR (x_counter >= 1488 AND x_counter <= 1505) OR (x_counter >= 1509 AND x_counter <= 1514) OR (x_counter >= 1518 AND x_counter <= 1523) OR (x_counter >= 1605 AND x_counter <= 1622) OR (x_counter >= 1626 AND x_counter <= 1631) OR (x_counter >= 1635 AND x_counter <= 1640)))
											OR	(y_counter = 364 AND ((x_counter >= 208 AND x_counter <= 225) OR (x_counter >= 229 AND x_counter <= 234) OR (x_counter >= 238 AND x_counter <= 243) OR (x_counter >= 325 AND x_counter <= 342) OR (x_counter >= 346 AND x_counter <= 351) OR (x_counter >= 355 AND x_counter <= 360) OR (x_counter >= 848 AND x_counter <= 865) OR (x_counter >= 869 AND x_counter <= 874) OR (x_counter >= 878 AND x_counter <= 883) OR (x_counter >= 965 AND x_counter <= 982) OR (x_counter >= 986 AND x_counter <= 991) OR (x_counter >= 995 AND x_counter <= 1000) OR (x_counter >= 1488 AND x_counter <= 1505) OR (x_counter >= 1509 AND x_counter <= 1514) OR (x_counter >= 1518 AND x_counter <= 1523) OR (x_counter >= 1605 AND x_counter <= 1622) OR (x_counter >= 1626 AND x_counter <= 1631) OR (x_counter >= 1635 AND x_counter <= 1640)))
											OR	(y_counter = 365 AND ((x_counter >= 208 AND x_counter <= 225) OR (x_counter >= 229 AND x_counter <= 234) OR (x_counter >= 238 AND x_counter <= 243) OR (x_counter >= 325 AND x_counter <= 342) OR (x_counter >= 346 AND x_counter <= 351) OR (x_counter >= 355 AND x_counter <= 360) OR (x_counter >= 848 AND x_counter <= 865) OR (x_counter >= 869 AND x_counter <= 874) OR (x_counter >= 878 AND x_counter <= 883) OR (x_counter >= 965 AND x_counter <= 982) OR (x_counter >= 986 AND x_counter <= 991) OR (x_counter >= 995 AND x_counter <= 1000) OR (x_counter >= 1488 AND x_counter <= 1505) OR (x_counter >= 1509 AND x_counter <= 1514) OR (x_counter >= 1518 AND x_counter <= 1523) OR (x_counter >= 1605 AND x_counter <= 1622) OR (x_counter >= 1626 AND x_counter <= 1631) OR (x_counter >= 1635 AND x_counter <= 1640)))
											OR	(y_counter = 366 AND ((x_counter >= 208 AND x_counter <= 225) OR (x_counter >= 229 AND x_counter <= 234) OR (x_counter >= 238 AND x_counter <= 243) OR (x_counter >= 325 AND x_counter <= 342) OR (x_counter >= 346 AND x_counter <= 351) OR (x_counter >= 355 AND x_counter <= 360) OR (x_counter >= 848 AND x_counter <= 865) OR (x_counter >= 869 AND x_counter <= 874) OR (x_counter >= 878 AND x_counter <= 883) OR (x_counter >= 965 AND x_counter <= 982) OR (x_counter >= 986 AND x_counter <= 991) OR (x_counter >= 995 AND x_counter <= 1000) OR (x_counter >= 1488 AND x_counter <= 1505) OR (x_counter >= 1509 AND x_counter <= 1514) OR (x_counter >= 1518 AND x_counter <= 1523) OR (x_counter >= 1605 AND x_counter <= 1622) OR (x_counter >= 1626 AND x_counter <= 1631) OR (x_counter >= 1635 AND x_counter <= 1640)))
											OR	(y_counter = 367 AND ((x_counter >= 208 AND x_counter <= 225) OR (x_counter >= 229 AND x_counter <= 234) OR (x_counter >= 238 AND x_counter <= 243) OR (x_counter >= 325 AND x_counter <= 342) OR (x_counter >= 346 AND x_counter <= 351) OR (x_counter >= 355 AND x_counter <= 360) OR (x_counter >= 848 AND x_counter <= 865) OR (x_counter >= 869 AND x_counter <= 874) OR (x_counter >= 878 AND x_counter <= 883) OR (x_counter >= 965 AND x_counter <= 982) OR (x_counter >= 986 AND x_counter <= 991) OR (x_counter >= 995 AND x_counter <= 1000) OR (x_counter >= 1488 AND x_counter <= 1505) OR (x_counter >= 1509 AND x_counter <= 1514) OR (x_counter >= 1518 AND x_counter <= 1523) OR (x_counter >= 1605 AND x_counter <= 1622) OR (x_counter >= 1626 AND x_counter <= 1631) OR (x_counter >= 1635 AND x_counter <= 1640)))
											OR	(y_counter = 368 AND ((x_counter >= 208 AND x_counter <= 213) OR (x_counter >= 220 AND x_counter <= 225) OR (x_counter >= 229 AND x_counter <= 234) OR (x_counter >= 325 AND x_counter <= 330) OR (x_counter >= 337 AND x_counter <= 342) OR (x_counter >= 346 AND x_counter <= 351) OR (x_counter >= 848 AND x_counter <= 853) OR (x_counter >= 860 AND x_counter <= 865) OR (x_counter >= 869 AND x_counter <= 874) OR (x_counter >= 965 AND x_counter <= 970) OR (x_counter >= 977 AND x_counter <= 982) OR (x_counter >= 986 AND x_counter <= 991) OR (x_counter >= 1488 AND x_counter <= 1493) OR (x_counter >= 1500 AND x_counter <= 1505) OR (x_counter >= 1509 AND x_counter <= 1514) OR (x_counter >= 1605 AND x_counter <= 1610) OR (x_counter >= 1617 AND x_counter <= 1622) OR (x_counter >= 1626 AND x_counter <= 1631)))
											OR	(y_counter = 369 AND ((x_counter >= 208 AND x_counter <= 213) OR (x_counter >= 220 AND x_counter <= 225) OR (x_counter >= 229 AND x_counter <= 234) OR (x_counter >= 325 AND x_counter <= 330) OR (x_counter >= 337 AND x_counter <= 342) OR (x_counter >= 346 AND x_counter <= 351) OR (x_counter >= 848 AND x_counter <= 853) OR (x_counter >= 860 AND x_counter <= 865) OR (x_counter >= 869 AND x_counter <= 874) OR (x_counter >= 965 AND x_counter <= 970) OR (x_counter >= 977 AND x_counter <= 982) OR (x_counter >= 986 AND x_counter <= 991) OR (x_counter >= 1488 AND x_counter <= 1493) OR (x_counter >= 1500 AND x_counter <= 1505) OR (x_counter >= 1509 AND x_counter <= 1514) OR (x_counter >= 1605 AND x_counter <= 1610) OR (x_counter >= 1617 AND x_counter <= 1622) OR (x_counter >= 1626 AND x_counter <= 1631)))
											OR	(y_counter = 370 AND ((x_counter >= 208 AND x_counter <= 213) OR (x_counter >= 220 AND x_counter <= 225) OR (x_counter >= 229 AND x_counter <= 234) OR (x_counter >= 325 AND x_counter <= 330) OR (x_counter >= 337 AND x_counter <= 342) OR (x_counter >= 346 AND x_counter <= 351) OR (x_counter >= 848 AND x_counter <= 853) OR (x_counter >= 860 AND x_counter <= 865) OR (x_counter >= 869 AND x_counter <= 874) OR (x_counter >= 965 AND x_counter <= 970) OR (x_counter >= 977 AND x_counter <= 982) OR (x_counter >= 986 AND x_counter <= 991) OR (x_counter >= 1488 AND x_counter <= 1493) OR (x_counter >= 1500 AND x_counter <= 1505) OR (x_counter >= 1509 AND x_counter <= 1514) OR (x_counter >= 1605 AND x_counter <= 1610) OR (x_counter >= 1617 AND x_counter <= 1622) OR (x_counter >= 1626 AND x_counter <= 1631)))
											OR	(y_counter = 371 AND ((x_counter >= 208 AND x_counter <= 213) OR (x_counter >= 220 AND x_counter <= 225) OR (x_counter >= 229 AND x_counter <= 234) OR (x_counter >= 238 AND x_counter <= 243) OR (x_counter >= 247 AND x_counter <= 258) OR (x_counter >= 262 AND x_counter <= 276) OR (x_counter >= 280 AND x_counter <= 294) OR (x_counter >= 298 AND x_counter <= 312) OR (x_counter >= 325 AND x_counter <= 330) OR (x_counter >= 337 AND x_counter <= 342) OR (x_counter >= 346 AND x_counter <= 351) OR (x_counter >= 355 AND x_counter <= 360) OR (x_counter >= 364 AND x_counter <= 378) OR (x_counter >= 382 AND x_counter <= 396) OR (x_counter >= 400 AND x_counter <= 405) OR (x_counter >= 409 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 429) OR (x_counter >= 848 AND x_counter <= 853) OR (x_counter >= 860 AND x_counter <= 865) OR (x_counter >= 869 AND x_counter <= 874) OR (x_counter >= 878 AND x_counter <= 883) OR (x_counter >= 887 AND x_counter <= 898) OR (x_counter >= 902 AND x_counter <= 916) OR (x_counter >= 920 AND x_counter <= 934) OR (x_counter >= 938 AND x_counter <= 952) OR (x_counter >= 965 AND x_counter <= 970) OR (x_counter >= 977 AND x_counter <= 982) OR (x_counter >= 986 AND x_counter <= 991) OR (x_counter >= 995 AND x_counter <= 1000) OR (x_counter >= 1004 AND x_counter <= 1018) OR (x_counter >= 1022 AND x_counter <= 1036) OR (x_counter >= 1040 AND x_counter <= 1045) OR (x_counter >= 1049 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1069) OR (x_counter >= 1488 AND x_counter <= 1493) OR (x_counter >= 1500 AND x_counter <= 1505) OR (x_counter >= 1509 AND x_counter <= 1514) OR (x_counter >= 1518 AND x_counter <= 1523) OR (x_counter >= 1527 AND x_counter <= 1538) OR (x_counter >= 1542 AND x_counter <= 1556) OR (x_counter >= 1560 AND x_counter <= 1574) OR (x_counter >= 1578 AND x_counter <= 1592) OR (x_counter >= 1605 AND x_counter <= 1610) OR (x_counter >= 1617 AND x_counter <= 1622) OR (x_counter >= 1626 AND x_counter <= 1631) OR (x_counter >= 1635 AND x_counter <= 1640) OR (x_counter >= 1644 AND x_counter <= 1658) OR (x_counter >= 1662 AND x_counter <= 1676) OR (x_counter >= 1680 AND x_counter <= 1685) OR (x_counter >= 1689 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1709)))
											OR	(y_counter = 372 AND ((x_counter >= 208 AND x_counter <= 213) OR (x_counter >= 220 AND x_counter <= 225) OR (x_counter >= 229 AND x_counter <= 234) OR (x_counter >= 238 AND x_counter <= 243) OR (x_counter >= 247 AND x_counter <= 258) OR (x_counter >= 262 AND x_counter <= 276) OR (x_counter >= 280 AND x_counter <= 294) OR (x_counter >= 298 AND x_counter <= 312) OR (x_counter >= 325 AND x_counter <= 330) OR (x_counter >= 337 AND x_counter <= 342) OR (x_counter >= 346 AND x_counter <= 351) OR (x_counter >= 355 AND x_counter <= 360) OR (x_counter >= 364 AND x_counter <= 378) OR (x_counter >= 382 AND x_counter <= 396) OR (x_counter >= 400 AND x_counter <= 405) OR (x_counter >= 409 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 429) OR (x_counter >= 848 AND x_counter <= 853) OR (x_counter >= 860 AND x_counter <= 865) OR (x_counter >= 869 AND x_counter <= 874) OR (x_counter >= 878 AND x_counter <= 883) OR (x_counter >= 887 AND x_counter <= 898) OR (x_counter >= 902 AND x_counter <= 916) OR (x_counter >= 920 AND x_counter <= 934) OR (x_counter >= 938 AND x_counter <= 952) OR (x_counter >= 965 AND x_counter <= 970) OR (x_counter >= 977 AND x_counter <= 982) OR (x_counter >= 986 AND x_counter <= 991) OR (x_counter >= 995 AND x_counter <= 1000) OR (x_counter >= 1004 AND x_counter <= 1018) OR (x_counter >= 1022 AND x_counter <= 1036) OR (x_counter >= 1040 AND x_counter <= 1045) OR (x_counter >= 1049 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1069) OR (x_counter >= 1488 AND x_counter <= 1493) OR (x_counter >= 1500 AND x_counter <= 1505) OR (x_counter >= 1509 AND x_counter <= 1514) OR (x_counter >= 1518 AND x_counter <= 1523) OR (x_counter >= 1527 AND x_counter <= 1538) OR (x_counter >= 1542 AND x_counter <= 1556) OR (x_counter >= 1560 AND x_counter <= 1574) OR (x_counter >= 1578 AND x_counter <= 1592) OR (x_counter >= 1605 AND x_counter <= 1610) OR (x_counter >= 1617 AND x_counter <= 1622) OR (x_counter >= 1626 AND x_counter <= 1631) OR (x_counter >= 1635 AND x_counter <= 1640) OR (x_counter >= 1644 AND x_counter <= 1658) OR (x_counter >= 1662 AND x_counter <= 1676) OR (x_counter >= 1680 AND x_counter <= 1685) OR (x_counter >= 1689 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1709)))
											OR	(y_counter = 373 AND ((x_counter >= 208 AND x_counter <= 213) OR (x_counter >= 220 AND x_counter <= 225) OR (x_counter >= 229 AND x_counter <= 234) OR (x_counter >= 238 AND x_counter <= 243) OR (x_counter >= 247 AND x_counter <= 258) OR (x_counter >= 262 AND x_counter <= 276) OR (x_counter >= 280 AND x_counter <= 294) OR (x_counter >= 298 AND x_counter <= 312) OR (x_counter >= 325 AND x_counter <= 330) OR (x_counter >= 337 AND x_counter <= 342) OR (x_counter >= 346 AND x_counter <= 351) OR (x_counter >= 355 AND x_counter <= 360) OR (x_counter >= 364 AND x_counter <= 378) OR (x_counter >= 382 AND x_counter <= 396) OR (x_counter >= 400 AND x_counter <= 405) OR (x_counter >= 409 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 429) OR (x_counter >= 848 AND x_counter <= 853) OR (x_counter >= 860 AND x_counter <= 865) OR (x_counter >= 869 AND x_counter <= 874) OR (x_counter >= 878 AND x_counter <= 883) OR (x_counter >= 887 AND x_counter <= 898) OR (x_counter >= 902 AND x_counter <= 916) OR (x_counter >= 920 AND x_counter <= 934) OR (x_counter >= 938 AND x_counter <= 952) OR (x_counter >= 965 AND x_counter <= 970) OR (x_counter >= 977 AND x_counter <= 982) OR (x_counter >= 986 AND x_counter <= 991) OR (x_counter >= 995 AND x_counter <= 1000) OR (x_counter >= 1004 AND x_counter <= 1018) OR (x_counter >= 1022 AND x_counter <= 1036) OR (x_counter >= 1040 AND x_counter <= 1045) OR (x_counter >= 1049 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1069) OR (x_counter >= 1488 AND x_counter <= 1493) OR (x_counter >= 1500 AND x_counter <= 1505) OR (x_counter >= 1509 AND x_counter <= 1514) OR (x_counter >= 1518 AND x_counter <= 1523) OR (x_counter >= 1527 AND x_counter <= 1538) OR (x_counter >= 1542 AND x_counter <= 1556) OR (x_counter >= 1560 AND x_counter <= 1574) OR (x_counter >= 1578 AND x_counter <= 1592) OR (x_counter >= 1605 AND x_counter <= 1610) OR (x_counter >= 1617 AND x_counter <= 1622) OR (x_counter >= 1626 AND x_counter <= 1631) OR (x_counter >= 1635 AND x_counter <= 1640) OR (x_counter >= 1644 AND x_counter <= 1658) OR (x_counter >= 1662 AND x_counter <= 1676) OR (x_counter >= 1680 AND x_counter <= 1685) OR (x_counter >= 1689 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1709)))
											OR	(y_counter = 374 AND ((x_counter >= 208 AND x_counter <= 225) OR (x_counter >= 229 AND x_counter <= 234) OR (x_counter >= 238 AND x_counter <= 243) OR (x_counter >= 247 AND x_counter <= 258) OR (x_counter >= 262 AND x_counter <= 276) OR (x_counter >= 280 AND x_counter <= 294) OR (x_counter >= 298 AND x_counter <= 312) OR (x_counter >= 325 AND x_counter <= 342) OR (x_counter >= 346 AND x_counter <= 351) OR (x_counter >= 355 AND x_counter <= 360) OR (x_counter >= 364 AND x_counter <= 378) OR (x_counter >= 382 AND x_counter <= 396) OR (x_counter >= 400 AND x_counter <= 405) OR (x_counter >= 409 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 429) OR (x_counter >= 848 AND x_counter <= 865) OR (x_counter >= 869 AND x_counter <= 874) OR (x_counter >= 878 AND x_counter <= 883) OR (x_counter >= 887 AND x_counter <= 898) OR (x_counter >= 902 AND x_counter <= 916) OR (x_counter >= 920 AND x_counter <= 934) OR (x_counter >= 938 AND x_counter <= 952) OR (x_counter >= 965 AND x_counter <= 982) OR (x_counter >= 986 AND x_counter <= 991) OR (x_counter >= 995 AND x_counter <= 1000) OR (x_counter >= 1004 AND x_counter <= 1018) OR (x_counter >= 1022 AND x_counter <= 1036) OR (x_counter >= 1040 AND x_counter <= 1045) OR (x_counter >= 1049 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1069) OR (x_counter >= 1488 AND x_counter <= 1505) OR (x_counter >= 1509 AND x_counter <= 1514) OR (x_counter >= 1518 AND x_counter <= 1523) OR (x_counter >= 1527 AND x_counter <= 1538) OR (x_counter >= 1542 AND x_counter <= 1556) OR (x_counter >= 1560 AND x_counter <= 1574) OR (x_counter >= 1578 AND x_counter <= 1592) OR (x_counter >= 1605 AND x_counter <= 1622) OR (x_counter >= 1626 AND x_counter <= 1631) OR (x_counter >= 1635 AND x_counter <= 1640) OR (x_counter >= 1644 AND x_counter <= 1658) OR (x_counter >= 1662 AND x_counter <= 1676) OR (x_counter >= 1680 AND x_counter <= 1685) OR (x_counter >= 1689 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1709)))
											OR	(y_counter = 375 AND ((x_counter >= 208 AND x_counter <= 225) OR (x_counter >= 229 AND x_counter <= 234) OR (x_counter >= 238 AND x_counter <= 243) OR (x_counter >= 247 AND x_counter <= 258) OR (x_counter >= 262 AND x_counter <= 276) OR (x_counter >= 280 AND x_counter <= 294) OR (x_counter >= 298 AND x_counter <= 312) OR (x_counter >= 325 AND x_counter <= 342) OR (x_counter >= 346 AND x_counter <= 351) OR (x_counter >= 355 AND x_counter <= 360) OR (x_counter >= 364 AND x_counter <= 378) OR (x_counter >= 382 AND x_counter <= 396) OR (x_counter >= 400 AND x_counter <= 405) OR (x_counter >= 409 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 429) OR (x_counter >= 848 AND x_counter <= 865) OR (x_counter >= 869 AND x_counter <= 874) OR (x_counter >= 878 AND x_counter <= 883) OR (x_counter >= 887 AND x_counter <= 898) OR (x_counter >= 902 AND x_counter <= 916) OR (x_counter >= 920 AND x_counter <= 934) OR (x_counter >= 938 AND x_counter <= 952) OR (x_counter >= 965 AND x_counter <= 982) OR (x_counter >= 986 AND x_counter <= 991) OR (x_counter >= 995 AND x_counter <= 1000) OR (x_counter >= 1004 AND x_counter <= 1018) OR (x_counter >= 1022 AND x_counter <= 1036) OR (x_counter >= 1040 AND x_counter <= 1045) OR (x_counter >= 1049 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1069) OR (x_counter >= 1488 AND x_counter <= 1505) OR (x_counter >= 1509 AND x_counter <= 1514) OR (x_counter >= 1518 AND x_counter <= 1523) OR (x_counter >= 1527 AND x_counter <= 1538) OR (x_counter >= 1542 AND x_counter <= 1556) OR (x_counter >= 1560 AND x_counter <= 1574) OR (x_counter >= 1578 AND x_counter <= 1592) OR (x_counter >= 1605 AND x_counter <= 1622) OR (x_counter >= 1626 AND x_counter <= 1631) OR (x_counter >= 1635 AND x_counter <= 1640) OR (x_counter >= 1644 AND x_counter <= 1658) OR (x_counter >= 1662 AND x_counter <= 1676) OR (x_counter >= 1680 AND x_counter <= 1685) OR (x_counter >= 1689 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1709)))
											OR	(y_counter = 376 AND ((x_counter >= 208 AND x_counter <= 225) OR (x_counter >= 229 AND x_counter <= 234) OR (x_counter >= 238 AND x_counter <= 243) OR (x_counter >= 247 AND x_counter <= 258) OR (x_counter >= 262 AND x_counter <= 276) OR (x_counter >= 280 AND x_counter <= 294) OR (x_counter >= 298 AND x_counter <= 312) OR (x_counter >= 325 AND x_counter <= 342) OR (x_counter >= 346 AND x_counter <= 351) OR (x_counter >= 355 AND x_counter <= 360) OR (x_counter >= 364 AND x_counter <= 378) OR (x_counter >= 382 AND x_counter <= 396) OR (x_counter >= 400 AND x_counter <= 405) OR (x_counter >= 409 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 429) OR (x_counter >= 848 AND x_counter <= 865) OR (x_counter >= 869 AND x_counter <= 874) OR (x_counter >= 878 AND x_counter <= 883) OR (x_counter >= 887 AND x_counter <= 898) OR (x_counter >= 902 AND x_counter <= 916) OR (x_counter >= 920 AND x_counter <= 934) OR (x_counter >= 938 AND x_counter <= 952) OR (x_counter >= 965 AND x_counter <= 982) OR (x_counter >= 986 AND x_counter <= 991) OR (x_counter >= 995 AND x_counter <= 1000) OR (x_counter >= 1004 AND x_counter <= 1018) OR (x_counter >= 1022 AND x_counter <= 1036) OR (x_counter >= 1040 AND x_counter <= 1045) OR (x_counter >= 1049 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1069) OR (x_counter >= 1488 AND x_counter <= 1505) OR (x_counter >= 1509 AND x_counter <= 1514) OR (x_counter >= 1518 AND x_counter <= 1523) OR (x_counter >= 1527 AND x_counter <= 1538) OR (x_counter >= 1542 AND x_counter <= 1556) OR (x_counter >= 1560 AND x_counter <= 1574) OR (x_counter >= 1578 AND x_counter <= 1592) OR (x_counter >= 1605 AND x_counter <= 1622) OR (x_counter >= 1626 AND x_counter <= 1631) OR (x_counter >= 1635 AND x_counter <= 1640) OR (x_counter >= 1644 AND x_counter <= 1658) OR (x_counter >= 1662 AND x_counter <= 1676) OR (x_counter >= 1680 AND x_counter <= 1685) OR (x_counter >= 1689 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1709)))
											OR	(y_counter = 377 AND ((x_counter >= 208 AND x_counter <= 225) OR (x_counter >= 229 AND x_counter <= 234) OR (x_counter >= 238 AND x_counter <= 243) OR (x_counter >= 247 AND x_counter <= 252) OR (x_counter >= 262 AND x_counter <= 267) OR (x_counter >= 271 AND x_counter <= 276) OR (x_counter >= 289 AND x_counter <= 294) OR (x_counter >= 307 AND x_counter <= 312) OR (x_counter >= 325 AND x_counter <= 342) OR (x_counter >= 346 AND x_counter <= 351) OR (x_counter >= 355 AND x_counter <= 360) OR (x_counter >= 364 AND x_counter <= 369) OR (x_counter >= 373 AND x_counter <= 378) OR (x_counter >= 382 AND x_counter <= 387) OR (x_counter >= 391 AND x_counter <= 396) OR (x_counter >= 400 AND x_counter <= 405) OR (x_counter >= 409 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 423) OR (x_counter >= 848 AND x_counter <= 865) OR (x_counter >= 869 AND x_counter <= 874) OR (x_counter >= 878 AND x_counter <= 883) OR (x_counter >= 887 AND x_counter <= 892) OR (x_counter >= 902 AND x_counter <= 907) OR (x_counter >= 911 AND x_counter <= 916) OR (x_counter >= 929 AND x_counter <= 934) OR (x_counter >= 947 AND x_counter <= 952) OR (x_counter >= 965 AND x_counter <= 982) OR (x_counter >= 986 AND x_counter <= 991) OR (x_counter >= 995 AND x_counter <= 1000) OR (x_counter >= 1004 AND x_counter <= 1009) OR (x_counter >= 1013 AND x_counter <= 1018) OR (x_counter >= 1022 AND x_counter <= 1027) OR (x_counter >= 1031 AND x_counter <= 1036) OR (x_counter >= 1040 AND x_counter <= 1045) OR (x_counter >= 1049 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1063) OR (x_counter >= 1488 AND x_counter <= 1505) OR (x_counter >= 1509 AND x_counter <= 1514) OR (x_counter >= 1518 AND x_counter <= 1523) OR (x_counter >= 1527 AND x_counter <= 1532) OR (x_counter >= 1542 AND x_counter <= 1547) OR (x_counter >= 1551 AND x_counter <= 1556) OR (x_counter >= 1569 AND x_counter <= 1574) OR (x_counter >= 1587 AND x_counter <= 1592) OR (x_counter >= 1605 AND x_counter <= 1622) OR (x_counter >= 1626 AND x_counter <= 1631) OR (x_counter >= 1635 AND x_counter <= 1640) OR (x_counter >= 1644 AND x_counter <= 1649) OR (x_counter >= 1653 AND x_counter <= 1658) OR (x_counter >= 1662 AND x_counter <= 1667) OR (x_counter >= 1671 AND x_counter <= 1676) OR (x_counter >= 1680 AND x_counter <= 1685) OR (x_counter >= 1689 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1703)))
											OR	(y_counter = 378 AND ((x_counter >= 208 AND x_counter <= 225) OR (x_counter >= 229 AND x_counter <= 234) OR (x_counter >= 238 AND x_counter <= 243) OR (x_counter >= 247 AND x_counter <= 252) OR (x_counter >= 262 AND x_counter <= 267) OR (x_counter >= 271 AND x_counter <= 276) OR (x_counter >= 289 AND x_counter <= 294) OR (x_counter >= 307 AND x_counter <= 312) OR (x_counter >= 325 AND x_counter <= 342) OR (x_counter >= 346 AND x_counter <= 351) OR (x_counter >= 355 AND x_counter <= 360) OR (x_counter >= 364 AND x_counter <= 369) OR (x_counter >= 373 AND x_counter <= 378) OR (x_counter >= 382 AND x_counter <= 387) OR (x_counter >= 391 AND x_counter <= 396) OR (x_counter >= 400 AND x_counter <= 405) OR (x_counter >= 409 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 423) OR (x_counter >= 848 AND x_counter <= 865) OR (x_counter >= 869 AND x_counter <= 874) OR (x_counter >= 878 AND x_counter <= 883) OR (x_counter >= 887 AND x_counter <= 892) OR (x_counter >= 902 AND x_counter <= 907) OR (x_counter >= 911 AND x_counter <= 916) OR (x_counter >= 929 AND x_counter <= 934) OR (x_counter >= 947 AND x_counter <= 952) OR (x_counter >= 965 AND x_counter <= 982) OR (x_counter >= 986 AND x_counter <= 991) OR (x_counter >= 995 AND x_counter <= 1000) OR (x_counter >= 1004 AND x_counter <= 1009) OR (x_counter >= 1013 AND x_counter <= 1018) OR (x_counter >= 1022 AND x_counter <= 1027) OR (x_counter >= 1031 AND x_counter <= 1036) OR (x_counter >= 1040 AND x_counter <= 1045) OR (x_counter >= 1049 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1063) OR (x_counter >= 1488 AND x_counter <= 1505) OR (x_counter >= 1509 AND x_counter <= 1514) OR (x_counter >= 1518 AND x_counter <= 1523) OR (x_counter >= 1527 AND x_counter <= 1532) OR (x_counter >= 1542 AND x_counter <= 1547) OR (x_counter >= 1551 AND x_counter <= 1556) OR (x_counter >= 1569 AND x_counter <= 1574) OR (x_counter >= 1587 AND x_counter <= 1592) OR (x_counter >= 1605 AND x_counter <= 1622) OR (x_counter >= 1626 AND x_counter <= 1631) OR (x_counter >= 1635 AND x_counter <= 1640) OR (x_counter >= 1644 AND x_counter <= 1649) OR (x_counter >= 1653 AND x_counter <= 1658) OR (x_counter >= 1662 AND x_counter <= 1667) OR (x_counter >= 1671 AND x_counter <= 1676) OR (x_counter >= 1680 AND x_counter <= 1685) OR (x_counter >= 1689 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1703)))
											OR	(y_counter = 379 AND ((x_counter >= 208 AND x_counter <= 225) OR (x_counter >= 229 AND x_counter <= 234) OR (x_counter >= 238 AND x_counter <= 243) OR (x_counter >= 247 AND x_counter <= 252) OR (x_counter >= 262 AND x_counter <= 267) OR (x_counter >= 271 AND x_counter <= 276) OR (x_counter >= 289 AND x_counter <= 294) OR (x_counter >= 307 AND x_counter <= 312) OR (x_counter >= 325 AND x_counter <= 342) OR (x_counter >= 346 AND x_counter <= 351) OR (x_counter >= 355 AND x_counter <= 360) OR (x_counter >= 364 AND x_counter <= 369) OR (x_counter >= 373 AND x_counter <= 378) OR (x_counter >= 382 AND x_counter <= 387) OR (x_counter >= 391 AND x_counter <= 396) OR (x_counter >= 400 AND x_counter <= 405) OR (x_counter >= 409 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 423) OR (x_counter >= 848 AND x_counter <= 865) OR (x_counter >= 869 AND x_counter <= 874) OR (x_counter >= 878 AND x_counter <= 883) OR (x_counter >= 887 AND x_counter <= 892) OR (x_counter >= 902 AND x_counter <= 907) OR (x_counter >= 911 AND x_counter <= 916) OR (x_counter >= 929 AND x_counter <= 934) OR (x_counter >= 947 AND x_counter <= 952) OR (x_counter >= 965 AND x_counter <= 982) OR (x_counter >= 986 AND x_counter <= 991) OR (x_counter >= 995 AND x_counter <= 1000) OR (x_counter >= 1004 AND x_counter <= 1009) OR (x_counter >= 1013 AND x_counter <= 1018) OR (x_counter >= 1022 AND x_counter <= 1027) OR (x_counter >= 1031 AND x_counter <= 1036) OR (x_counter >= 1040 AND x_counter <= 1045) OR (x_counter >= 1049 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1063) OR (x_counter >= 1488 AND x_counter <= 1505) OR (x_counter >= 1509 AND x_counter <= 1514) OR (x_counter >= 1518 AND x_counter <= 1523) OR (x_counter >= 1527 AND x_counter <= 1532) OR (x_counter >= 1542 AND x_counter <= 1547) OR (x_counter >= 1551 AND x_counter <= 1556) OR (x_counter >= 1569 AND x_counter <= 1574) OR (x_counter >= 1587 AND x_counter <= 1592) OR (x_counter >= 1605 AND x_counter <= 1622) OR (x_counter >= 1626 AND x_counter <= 1631) OR (x_counter >= 1635 AND x_counter <= 1640) OR (x_counter >= 1644 AND x_counter <= 1649) OR (x_counter >= 1653 AND x_counter <= 1658) OR (x_counter >= 1662 AND x_counter <= 1667) OR (x_counter >= 1671 AND x_counter <= 1676) OR (x_counter >= 1680 AND x_counter <= 1685) OR (x_counter >= 1689 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1703)))
											OR	(y_counter = 380 AND ((x_counter >= 208 AND x_counter <= 213) OR (x_counter >= 220 AND x_counter <= 225) OR (x_counter >= 229 AND x_counter <= 234) OR (x_counter >= 238 AND x_counter <= 243) OR (x_counter >= 247 AND x_counter <= 252) OR (x_counter >= 262 AND x_counter <= 276) OR (x_counter >= 280 AND x_counter <= 294) OR (x_counter >= 298 AND x_counter <= 312) OR (x_counter >= 325 AND x_counter <= 330) OR (x_counter >= 337 AND x_counter <= 342) OR (x_counter >= 346 AND x_counter <= 351) OR (x_counter >= 355 AND x_counter <= 360) OR (x_counter >= 364 AND x_counter <= 369) OR (x_counter >= 373 AND x_counter <= 378) OR (x_counter >= 382 AND x_counter <= 387) OR (x_counter >= 391 AND x_counter <= 396) OR (x_counter >= 400 AND x_counter <= 405) OR (x_counter >= 409 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 423) OR (x_counter >= 848 AND x_counter <= 853) OR (x_counter >= 860 AND x_counter <= 865) OR (x_counter >= 869 AND x_counter <= 874) OR (x_counter >= 878 AND x_counter <= 883) OR (x_counter >= 887 AND x_counter <= 892) OR (x_counter >= 902 AND x_counter <= 916) OR (x_counter >= 920 AND x_counter <= 934) OR (x_counter >= 938 AND x_counter <= 952) OR (x_counter >= 965 AND x_counter <= 970) OR (x_counter >= 977 AND x_counter <= 982) OR (x_counter >= 986 AND x_counter <= 991) OR (x_counter >= 995 AND x_counter <= 1000) OR (x_counter >= 1004 AND x_counter <= 1009) OR (x_counter >= 1013 AND x_counter <= 1018) OR (x_counter >= 1022 AND x_counter <= 1027) OR (x_counter >= 1031 AND x_counter <= 1036) OR (x_counter >= 1040 AND x_counter <= 1045) OR (x_counter >= 1049 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1063) OR (x_counter >= 1488 AND x_counter <= 1493) OR (x_counter >= 1500 AND x_counter <= 1505) OR (x_counter >= 1509 AND x_counter <= 1514) OR (x_counter >= 1518 AND x_counter <= 1523) OR (x_counter >= 1527 AND x_counter <= 1532) OR (x_counter >= 1542 AND x_counter <= 1556) OR (x_counter >= 1560 AND x_counter <= 1574) OR (x_counter >= 1578 AND x_counter <= 1592) OR (x_counter >= 1605 AND x_counter <= 1610) OR (x_counter >= 1617 AND x_counter <= 1622) OR (x_counter >= 1626 AND x_counter <= 1631) OR (x_counter >= 1635 AND x_counter <= 1640) OR (x_counter >= 1644 AND x_counter <= 1649) OR (x_counter >= 1653 AND x_counter <= 1658) OR (x_counter >= 1662 AND x_counter <= 1667) OR (x_counter >= 1671 AND x_counter <= 1676) OR (x_counter >= 1680 AND x_counter <= 1685) OR (x_counter >= 1689 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1703)))
											OR	(y_counter = 381 AND ((x_counter >= 208 AND x_counter <= 213) OR (x_counter >= 220 AND x_counter <= 225) OR (x_counter >= 229 AND x_counter <= 234) OR (x_counter >= 238 AND x_counter <= 243) OR (x_counter >= 247 AND x_counter <= 252) OR (x_counter >= 262 AND x_counter <= 276) OR (x_counter >= 280 AND x_counter <= 294) OR (x_counter >= 298 AND x_counter <= 312) OR (x_counter >= 325 AND x_counter <= 330) OR (x_counter >= 337 AND x_counter <= 342) OR (x_counter >= 346 AND x_counter <= 351) OR (x_counter >= 355 AND x_counter <= 360) OR (x_counter >= 364 AND x_counter <= 369) OR (x_counter >= 373 AND x_counter <= 378) OR (x_counter >= 382 AND x_counter <= 387) OR (x_counter >= 391 AND x_counter <= 396) OR (x_counter >= 400 AND x_counter <= 405) OR (x_counter >= 409 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 423) OR (x_counter >= 848 AND x_counter <= 853) OR (x_counter >= 860 AND x_counter <= 865) OR (x_counter >= 869 AND x_counter <= 874) OR (x_counter >= 878 AND x_counter <= 883) OR (x_counter >= 887 AND x_counter <= 892) OR (x_counter >= 902 AND x_counter <= 916) OR (x_counter >= 920 AND x_counter <= 934) OR (x_counter >= 938 AND x_counter <= 952) OR (x_counter >= 965 AND x_counter <= 970) OR (x_counter >= 977 AND x_counter <= 982) OR (x_counter >= 986 AND x_counter <= 991) OR (x_counter >= 995 AND x_counter <= 1000) OR (x_counter >= 1004 AND x_counter <= 1009) OR (x_counter >= 1013 AND x_counter <= 1018) OR (x_counter >= 1022 AND x_counter <= 1027) OR (x_counter >= 1031 AND x_counter <= 1036) OR (x_counter >= 1040 AND x_counter <= 1045) OR (x_counter >= 1049 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1063) OR (x_counter >= 1488 AND x_counter <= 1493) OR (x_counter >= 1500 AND x_counter <= 1505) OR (x_counter >= 1509 AND x_counter <= 1514) OR (x_counter >= 1518 AND x_counter <= 1523) OR (x_counter >= 1527 AND x_counter <= 1532) OR (x_counter >= 1542 AND x_counter <= 1556) OR (x_counter >= 1560 AND x_counter <= 1574) OR (x_counter >= 1578 AND x_counter <= 1592) OR (x_counter >= 1605 AND x_counter <= 1610) OR (x_counter >= 1617 AND x_counter <= 1622) OR (x_counter >= 1626 AND x_counter <= 1631) OR (x_counter >= 1635 AND x_counter <= 1640) OR (x_counter >= 1644 AND x_counter <= 1649) OR (x_counter >= 1653 AND x_counter <= 1658) OR (x_counter >= 1662 AND x_counter <= 1667) OR (x_counter >= 1671 AND x_counter <= 1676) OR (x_counter >= 1680 AND x_counter <= 1685) OR (x_counter >= 1689 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1703)))
											OR	(y_counter = 382 AND ((x_counter >= 208 AND x_counter <= 213) OR (x_counter >= 220 AND x_counter <= 225) OR (x_counter >= 229 AND x_counter <= 234) OR (x_counter >= 238 AND x_counter <= 243) OR (x_counter >= 247 AND x_counter <= 252) OR (x_counter >= 262 AND x_counter <= 276) OR (x_counter >= 280 AND x_counter <= 294) OR (x_counter >= 298 AND x_counter <= 312) OR (x_counter >= 325 AND x_counter <= 330) OR (x_counter >= 337 AND x_counter <= 342) OR (x_counter >= 346 AND x_counter <= 351) OR (x_counter >= 355 AND x_counter <= 360) OR (x_counter >= 364 AND x_counter <= 369) OR (x_counter >= 373 AND x_counter <= 378) OR (x_counter >= 382 AND x_counter <= 387) OR (x_counter >= 391 AND x_counter <= 396) OR (x_counter >= 400 AND x_counter <= 405) OR (x_counter >= 409 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 423) OR (x_counter >= 848 AND x_counter <= 853) OR (x_counter >= 860 AND x_counter <= 865) OR (x_counter >= 869 AND x_counter <= 874) OR (x_counter >= 878 AND x_counter <= 883) OR (x_counter >= 887 AND x_counter <= 892) OR (x_counter >= 902 AND x_counter <= 916) OR (x_counter >= 920 AND x_counter <= 934) OR (x_counter >= 938 AND x_counter <= 952) OR (x_counter >= 965 AND x_counter <= 970) OR (x_counter >= 977 AND x_counter <= 982) OR (x_counter >= 986 AND x_counter <= 991) OR (x_counter >= 995 AND x_counter <= 1000) OR (x_counter >= 1004 AND x_counter <= 1009) OR (x_counter >= 1013 AND x_counter <= 1018) OR (x_counter >= 1022 AND x_counter <= 1027) OR (x_counter >= 1031 AND x_counter <= 1036) OR (x_counter >= 1040 AND x_counter <= 1045) OR (x_counter >= 1049 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1063) OR (x_counter >= 1488 AND x_counter <= 1493) OR (x_counter >= 1500 AND x_counter <= 1505) OR (x_counter >= 1509 AND x_counter <= 1514) OR (x_counter >= 1518 AND x_counter <= 1523) OR (x_counter >= 1527 AND x_counter <= 1532) OR (x_counter >= 1542 AND x_counter <= 1556) OR (x_counter >= 1560 AND x_counter <= 1574) OR (x_counter >= 1578 AND x_counter <= 1592) OR (x_counter >= 1605 AND x_counter <= 1610) OR (x_counter >= 1617 AND x_counter <= 1622) OR (x_counter >= 1626 AND x_counter <= 1631) OR (x_counter >= 1635 AND x_counter <= 1640) OR (x_counter >= 1644 AND x_counter <= 1649) OR (x_counter >= 1653 AND x_counter <= 1658) OR (x_counter >= 1662 AND x_counter <= 1667) OR (x_counter >= 1671 AND x_counter <= 1676) OR (x_counter >= 1680 AND x_counter <= 1685) OR (x_counter >= 1689 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1703)))
											OR	(y_counter = 383 AND ((x_counter >= 208 AND x_counter <= 213) OR (x_counter >= 220 AND x_counter <= 225) OR (x_counter >= 229 AND x_counter <= 234) OR (x_counter >= 238 AND x_counter <= 243) OR (x_counter >= 247 AND x_counter <= 252) OR (x_counter >= 262 AND x_counter <= 267) OR (x_counter >= 280 AND x_counter <= 285) OR (x_counter >= 298 AND x_counter <= 303) OR (x_counter >= 307 AND x_counter <= 312) OR (x_counter >= 325 AND x_counter <= 330) OR (x_counter >= 337 AND x_counter <= 342) OR (x_counter >= 346 AND x_counter <= 351) OR (x_counter >= 355 AND x_counter <= 360) OR (x_counter >= 364 AND x_counter <= 369) OR (x_counter >= 373 AND x_counter <= 378) OR (x_counter >= 382 AND x_counter <= 387) OR (x_counter >= 391 AND x_counter <= 396) OR (x_counter >= 400 AND x_counter <= 405) OR (x_counter >= 409 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 423) OR (x_counter >= 848 AND x_counter <= 853) OR (x_counter >= 860 AND x_counter <= 865) OR (x_counter >= 869 AND x_counter <= 874) OR (x_counter >= 878 AND x_counter <= 883) OR (x_counter >= 887 AND x_counter <= 892) OR (x_counter >= 902 AND x_counter <= 907) OR (x_counter >= 920 AND x_counter <= 925) OR (x_counter >= 938 AND x_counter <= 943) OR (x_counter >= 947 AND x_counter <= 952) OR (x_counter >= 965 AND x_counter <= 970) OR (x_counter >= 977 AND x_counter <= 982) OR (x_counter >= 986 AND x_counter <= 991) OR (x_counter >= 995 AND x_counter <= 1000) OR (x_counter >= 1004 AND x_counter <= 1009) OR (x_counter >= 1013 AND x_counter <= 1018) OR (x_counter >= 1022 AND x_counter <= 1027) OR (x_counter >= 1031 AND x_counter <= 1036) OR (x_counter >= 1040 AND x_counter <= 1045) OR (x_counter >= 1049 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1063) OR (x_counter >= 1488 AND x_counter <= 1493) OR (x_counter >= 1500 AND x_counter <= 1505) OR (x_counter >= 1509 AND x_counter <= 1514) OR (x_counter >= 1518 AND x_counter <= 1523) OR (x_counter >= 1527 AND x_counter <= 1532) OR (x_counter >= 1542 AND x_counter <= 1547) OR (x_counter >= 1560 AND x_counter <= 1565) OR (x_counter >= 1578 AND x_counter <= 1583) OR (x_counter >= 1587 AND x_counter <= 1592) OR (x_counter >= 1605 AND x_counter <= 1610) OR (x_counter >= 1617 AND x_counter <= 1622) OR (x_counter >= 1626 AND x_counter <= 1631) OR (x_counter >= 1635 AND x_counter <= 1640) OR (x_counter >= 1644 AND x_counter <= 1649) OR (x_counter >= 1653 AND x_counter <= 1658) OR (x_counter >= 1662 AND x_counter <= 1667) OR (x_counter >= 1671 AND x_counter <= 1676) OR (x_counter >= 1680 AND x_counter <= 1685) OR (x_counter >= 1689 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1703)))
											OR	(y_counter = 384 AND ((x_counter >= 208 AND x_counter <= 213) OR (x_counter >= 220 AND x_counter <= 225) OR (x_counter >= 229 AND x_counter <= 234) OR (x_counter >= 238 AND x_counter <= 243) OR (x_counter >= 247 AND x_counter <= 252) OR (x_counter >= 262 AND x_counter <= 267) OR (x_counter >= 280 AND x_counter <= 285) OR (x_counter >= 298 AND x_counter <= 303) OR (x_counter >= 307 AND x_counter <= 312) OR (x_counter >= 325 AND x_counter <= 330) OR (x_counter >= 337 AND x_counter <= 342) OR (x_counter >= 346 AND x_counter <= 351) OR (x_counter >= 355 AND x_counter <= 360) OR (x_counter >= 364 AND x_counter <= 369) OR (x_counter >= 373 AND x_counter <= 378) OR (x_counter >= 382 AND x_counter <= 387) OR (x_counter >= 391 AND x_counter <= 396) OR (x_counter >= 400 AND x_counter <= 405) OR (x_counter >= 409 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 423) OR (x_counter >= 848 AND x_counter <= 853) OR (x_counter >= 860 AND x_counter <= 865) OR (x_counter >= 869 AND x_counter <= 874) OR (x_counter >= 878 AND x_counter <= 883) OR (x_counter >= 887 AND x_counter <= 892) OR (x_counter >= 902 AND x_counter <= 907) OR (x_counter >= 920 AND x_counter <= 925) OR (x_counter >= 938 AND x_counter <= 943) OR (x_counter >= 947 AND x_counter <= 952) OR (x_counter >= 965 AND x_counter <= 970) OR (x_counter >= 977 AND x_counter <= 982) OR (x_counter >= 986 AND x_counter <= 991) OR (x_counter >= 995 AND x_counter <= 1000) OR (x_counter >= 1004 AND x_counter <= 1009) OR (x_counter >= 1013 AND x_counter <= 1018) OR (x_counter >= 1022 AND x_counter <= 1027) OR (x_counter >= 1031 AND x_counter <= 1036) OR (x_counter >= 1040 AND x_counter <= 1045) OR (x_counter >= 1049 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1063) OR (x_counter >= 1488 AND x_counter <= 1493) OR (x_counter >= 1500 AND x_counter <= 1505) OR (x_counter >= 1509 AND x_counter <= 1514) OR (x_counter >= 1518 AND x_counter <= 1523) OR (x_counter >= 1527 AND x_counter <= 1532) OR (x_counter >= 1542 AND x_counter <= 1547) OR (x_counter >= 1560 AND x_counter <= 1565) OR (x_counter >= 1578 AND x_counter <= 1583) OR (x_counter >= 1587 AND x_counter <= 1592) OR (x_counter >= 1605 AND x_counter <= 1610) OR (x_counter >= 1617 AND x_counter <= 1622) OR (x_counter >= 1626 AND x_counter <= 1631) OR (x_counter >= 1635 AND x_counter <= 1640) OR (x_counter >= 1644 AND x_counter <= 1649) OR (x_counter >= 1653 AND x_counter <= 1658) OR (x_counter >= 1662 AND x_counter <= 1667) OR (x_counter >= 1671 AND x_counter <= 1676) OR (x_counter >= 1680 AND x_counter <= 1685) OR (x_counter >= 1689 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1703)))
											OR	(y_counter = 385 AND ((x_counter >= 208 AND x_counter <= 213) OR (x_counter >= 220 AND x_counter <= 225) OR (x_counter >= 229 AND x_counter <= 234) OR (x_counter >= 238 AND x_counter <= 243) OR (x_counter >= 247 AND x_counter <= 252) OR (x_counter >= 262 AND x_counter <= 267) OR (x_counter >= 280 AND x_counter <= 285) OR (x_counter >= 298 AND x_counter <= 303) OR (x_counter >= 307 AND x_counter <= 312) OR (x_counter >= 325 AND x_counter <= 330) OR (x_counter >= 337 AND x_counter <= 342) OR (x_counter >= 346 AND x_counter <= 351) OR (x_counter >= 355 AND x_counter <= 360) OR (x_counter >= 364 AND x_counter <= 369) OR (x_counter >= 373 AND x_counter <= 378) OR (x_counter >= 382 AND x_counter <= 387) OR (x_counter >= 391 AND x_counter <= 396) OR (x_counter >= 400 AND x_counter <= 405) OR (x_counter >= 409 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 423) OR (x_counter >= 848 AND x_counter <= 853) OR (x_counter >= 860 AND x_counter <= 865) OR (x_counter >= 869 AND x_counter <= 874) OR (x_counter >= 878 AND x_counter <= 883) OR (x_counter >= 887 AND x_counter <= 892) OR (x_counter >= 902 AND x_counter <= 907) OR (x_counter >= 920 AND x_counter <= 925) OR (x_counter >= 938 AND x_counter <= 943) OR (x_counter >= 947 AND x_counter <= 952) OR (x_counter >= 965 AND x_counter <= 970) OR (x_counter >= 977 AND x_counter <= 982) OR (x_counter >= 986 AND x_counter <= 991) OR (x_counter >= 995 AND x_counter <= 1000) OR (x_counter >= 1004 AND x_counter <= 1009) OR (x_counter >= 1013 AND x_counter <= 1018) OR (x_counter >= 1022 AND x_counter <= 1027) OR (x_counter >= 1031 AND x_counter <= 1036) OR (x_counter >= 1040 AND x_counter <= 1045) OR (x_counter >= 1049 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1063) OR (x_counter >= 1488 AND x_counter <= 1493) OR (x_counter >= 1500 AND x_counter <= 1505) OR (x_counter >= 1509 AND x_counter <= 1514) OR (x_counter >= 1518 AND x_counter <= 1523) OR (x_counter >= 1527 AND x_counter <= 1532) OR (x_counter >= 1542 AND x_counter <= 1547) OR (x_counter >= 1560 AND x_counter <= 1565) OR (x_counter >= 1578 AND x_counter <= 1583) OR (x_counter >= 1587 AND x_counter <= 1592) OR (x_counter >= 1605 AND x_counter <= 1610) OR (x_counter >= 1617 AND x_counter <= 1622) OR (x_counter >= 1626 AND x_counter <= 1631) OR (x_counter >= 1635 AND x_counter <= 1640) OR (x_counter >= 1644 AND x_counter <= 1649) OR (x_counter >= 1653 AND x_counter <= 1658) OR (x_counter >= 1662 AND x_counter <= 1667) OR (x_counter >= 1671 AND x_counter <= 1676) OR (x_counter >= 1680 AND x_counter <= 1685) OR (x_counter >= 1689 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1703)))
											OR	(y_counter = 386 AND ((x_counter >= 208 AND x_counter <= 213) OR (x_counter >= 220 AND x_counter <= 225) OR (x_counter >= 229 AND x_counter <= 234) OR (x_counter >= 238 AND x_counter <= 243) OR (x_counter >= 247 AND x_counter <= 252) OR (x_counter >= 262 AND x_counter <= 276) OR (x_counter >= 280 AND x_counter <= 294) OR (x_counter >= 298 AND x_counter <= 312) OR (x_counter >= 325 AND x_counter <= 330) OR (x_counter >= 337 AND x_counter <= 342) OR (x_counter >= 346 AND x_counter <= 351) OR (x_counter >= 355 AND x_counter <= 360) OR (x_counter >= 364 AND x_counter <= 378) OR (x_counter >= 382 AND x_counter <= 396) OR (x_counter >= 400 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 423) OR (x_counter >= 848 AND x_counter <= 853) OR (x_counter >= 860 AND x_counter <= 865) OR (x_counter >= 869 AND x_counter <= 874) OR (x_counter >= 878 AND x_counter <= 883) OR (x_counter >= 887 AND x_counter <= 892) OR (x_counter >= 902 AND x_counter <= 916) OR (x_counter >= 920 AND x_counter <= 934) OR (x_counter >= 938 AND x_counter <= 952) OR (x_counter >= 965 AND x_counter <= 970) OR (x_counter >= 977 AND x_counter <= 982) OR (x_counter >= 986 AND x_counter <= 991) OR (x_counter >= 995 AND x_counter <= 1000) OR (x_counter >= 1004 AND x_counter <= 1018) OR (x_counter >= 1022 AND x_counter <= 1036) OR (x_counter >= 1040 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1063) OR (x_counter >= 1488 AND x_counter <= 1493) OR (x_counter >= 1500 AND x_counter <= 1505) OR (x_counter >= 1509 AND x_counter <= 1514) OR (x_counter >= 1518 AND x_counter <= 1523) OR (x_counter >= 1527 AND x_counter <= 1532) OR (x_counter >= 1542 AND x_counter <= 1556) OR (x_counter >= 1560 AND x_counter <= 1574) OR (x_counter >= 1578 AND x_counter <= 1592) OR (x_counter >= 1605 AND x_counter <= 1610) OR (x_counter >= 1617 AND x_counter <= 1622) OR (x_counter >= 1626 AND x_counter <= 1631) OR (x_counter >= 1635 AND x_counter <= 1640) OR (x_counter >= 1644 AND x_counter <= 1658) OR (x_counter >= 1662 AND x_counter <= 1676) OR (x_counter >= 1680 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1703)))
											OR	(y_counter = 387 AND ((x_counter >= 208 AND x_counter <= 213) OR (x_counter >= 220 AND x_counter <= 225) OR (x_counter >= 229 AND x_counter <= 234) OR (x_counter >= 238 AND x_counter <= 243) OR (x_counter >= 247 AND x_counter <= 252) OR (x_counter >= 262 AND x_counter <= 276) OR (x_counter >= 280 AND x_counter <= 294) OR (x_counter >= 298 AND x_counter <= 312) OR (x_counter >= 325 AND x_counter <= 330) OR (x_counter >= 337 AND x_counter <= 342) OR (x_counter >= 346 AND x_counter <= 351) OR (x_counter >= 355 AND x_counter <= 360) OR (x_counter >= 364 AND x_counter <= 378) OR (x_counter >= 382 AND x_counter <= 396) OR (x_counter >= 400 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 423) OR (x_counter >= 848 AND x_counter <= 853) OR (x_counter >= 860 AND x_counter <= 865) OR (x_counter >= 869 AND x_counter <= 874) OR (x_counter >= 878 AND x_counter <= 883) OR (x_counter >= 887 AND x_counter <= 892) OR (x_counter >= 902 AND x_counter <= 916) OR (x_counter >= 920 AND x_counter <= 934) OR (x_counter >= 938 AND x_counter <= 952) OR (x_counter >= 965 AND x_counter <= 970) OR (x_counter >= 977 AND x_counter <= 982) OR (x_counter >= 986 AND x_counter <= 991) OR (x_counter >= 995 AND x_counter <= 1000) OR (x_counter >= 1004 AND x_counter <= 1018) OR (x_counter >= 1022 AND x_counter <= 1036) OR (x_counter >= 1040 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1063) OR (x_counter >= 1488 AND x_counter <= 1493) OR (x_counter >= 1500 AND x_counter <= 1505) OR (x_counter >= 1509 AND x_counter <= 1514) OR (x_counter >= 1518 AND x_counter <= 1523) OR (x_counter >= 1527 AND x_counter <= 1532) OR (x_counter >= 1542 AND x_counter <= 1556) OR (x_counter >= 1560 AND x_counter <= 1574) OR (x_counter >= 1578 AND x_counter <= 1592) OR (x_counter >= 1605 AND x_counter <= 1610) OR (x_counter >= 1617 AND x_counter <= 1622) OR (x_counter >= 1626 AND x_counter <= 1631) OR (x_counter >= 1635 AND x_counter <= 1640) OR (x_counter >= 1644 AND x_counter <= 1658) OR (x_counter >= 1662 AND x_counter <= 1676) OR (x_counter >= 1680 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1703)))
											OR	(y_counter = 388 AND ((x_counter >= 208 AND x_counter <= 213) OR (x_counter >= 220 AND x_counter <= 225) OR (x_counter >= 229 AND x_counter <= 234) OR (x_counter >= 238 AND x_counter <= 243) OR (x_counter >= 247 AND x_counter <= 252) OR (x_counter >= 262 AND x_counter <= 276) OR (x_counter >= 280 AND x_counter <= 294) OR (x_counter >= 298 AND x_counter <= 312) OR (x_counter >= 325 AND x_counter <= 330) OR (x_counter >= 337 AND x_counter <= 342) OR (x_counter >= 346 AND x_counter <= 351) OR (x_counter >= 355 AND x_counter <= 360) OR (x_counter >= 364 AND x_counter <= 378) OR (x_counter >= 382 AND x_counter <= 396) OR (x_counter >= 400 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 423) OR (x_counter >= 848 AND x_counter <= 853) OR (x_counter >= 860 AND x_counter <= 865) OR (x_counter >= 869 AND x_counter <= 874) OR (x_counter >= 878 AND x_counter <= 883) OR (x_counter >= 887 AND x_counter <= 892) OR (x_counter >= 902 AND x_counter <= 916) OR (x_counter >= 920 AND x_counter <= 934) OR (x_counter >= 938 AND x_counter <= 952) OR (x_counter >= 965 AND x_counter <= 970) OR (x_counter >= 977 AND x_counter <= 982) OR (x_counter >= 986 AND x_counter <= 991) OR (x_counter >= 995 AND x_counter <= 1000) OR (x_counter >= 1004 AND x_counter <= 1018) OR (x_counter >= 1022 AND x_counter <= 1036) OR (x_counter >= 1040 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1063) OR (x_counter >= 1488 AND x_counter <= 1493) OR (x_counter >= 1500 AND x_counter <= 1505) OR (x_counter >= 1509 AND x_counter <= 1514) OR (x_counter >= 1518 AND x_counter <= 1523) OR (x_counter >= 1527 AND x_counter <= 1532) OR (x_counter >= 1542 AND x_counter <= 1556) OR (x_counter >= 1560 AND x_counter <= 1574) OR (x_counter >= 1578 AND x_counter <= 1592) OR (x_counter >= 1605 AND x_counter <= 1610) OR (x_counter >= 1617 AND x_counter <= 1622) OR (x_counter >= 1626 AND x_counter <= 1631) OR (x_counter >= 1635 AND x_counter <= 1640) OR (x_counter >= 1644 AND x_counter <= 1658) OR (x_counter >= 1662 AND x_counter <= 1676) OR (x_counter >= 1680 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1703)))
											OR	(y_counter = 389 AND ((x_counter >= 208 AND x_counter <= 213) OR (x_counter >= 220 AND x_counter <= 225) OR (x_counter >= 229 AND x_counter <= 234) OR (x_counter >= 238 AND x_counter <= 243) OR (x_counter >= 247 AND x_counter <= 252) OR (x_counter >= 262 AND x_counter <= 276) OR (x_counter >= 280 AND x_counter <= 294) OR (x_counter >= 298 AND x_counter <= 312) OR (x_counter >= 325 AND x_counter <= 330) OR (x_counter >= 337 AND x_counter <= 342) OR (x_counter >= 346 AND x_counter <= 351) OR (x_counter >= 355 AND x_counter <= 360) OR (x_counter >= 364 AND x_counter <= 378) OR (x_counter >= 382 AND x_counter <= 396) OR (x_counter >= 400 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 423) OR (x_counter >= 848 AND x_counter <= 853) OR (x_counter >= 860 AND x_counter <= 865) OR (x_counter >= 869 AND x_counter <= 874) OR (x_counter >= 878 AND x_counter <= 883) OR (x_counter >= 887 AND x_counter <= 892) OR (x_counter >= 902 AND x_counter <= 916) OR (x_counter >= 920 AND x_counter <= 934) OR (x_counter >= 938 AND x_counter <= 952) OR (x_counter >= 965 AND x_counter <= 970) OR (x_counter >= 977 AND x_counter <= 982) OR (x_counter >= 986 AND x_counter <= 991) OR (x_counter >= 995 AND x_counter <= 1000) OR (x_counter >= 1004 AND x_counter <= 1018) OR (x_counter >= 1022 AND x_counter <= 1036) OR (x_counter >= 1040 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1063) OR (x_counter >= 1488 AND x_counter <= 1493) OR (x_counter >= 1500 AND x_counter <= 1505) OR (x_counter >= 1509 AND x_counter <= 1514) OR (x_counter >= 1518 AND x_counter <= 1523) OR (x_counter >= 1527 AND x_counter <= 1532) OR (x_counter >= 1542 AND x_counter <= 1556) OR (x_counter >= 1560 AND x_counter <= 1574) OR (x_counter >= 1578 AND x_counter <= 1592) OR (x_counter >= 1605 AND x_counter <= 1610) OR (x_counter >= 1617 AND x_counter <= 1622) OR (x_counter >= 1626 AND x_counter <= 1631) OR (x_counter >= 1635 AND x_counter <= 1640) OR (x_counter >= 1644 AND x_counter <= 1658) OR (x_counter >= 1662 AND x_counter <= 1676) OR (x_counter >= 1680 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1703)))
											OR	(y_counter = 390 AND ((x_counter >= 208 AND x_counter <= 213) OR (x_counter >= 220 AND x_counter <= 225) OR (x_counter >= 229 AND x_counter <= 234) OR (x_counter >= 238 AND x_counter <= 243) OR (x_counter >= 247 AND x_counter <= 252) OR (x_counter >= 262 AND x_counter <= 276) OR (x_counter >= 280 AND x_counter <= 294) OR (x_counter >= 298 AND x_counter <= 312) OR (x_counter >= 325 AND x_counter <= 330) OR (x_counter >= 337 AND x_counter <= 342) OR (x_counter >= 346 AND x_counter <= 351) OR (x_counter >= 355 AND x_counter <= 360) OR (x_counter >= 364 AND x_counter <= 378) OR (x_counter >= 382 AND x_counter <= 396) OR (x_counter >= 400 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 423) OR (x_counter >= 848 AND x_counter <= 853) OR (x_counter >= 860 AND x_counter <= 865) OR (x_counter >= 869 AND x_counter <= 874) OR (x_counter >= 878 AND x_counter <= 883) OR (x_counter >= 887 AND x_counter <= 892) OR (x_counter >= 902 AND x_counter <= 916) OR (x_counter >= 920 AND x_counter <= 934) OR (x_counter >= 938 AND x_counter <= 952) OR (x_counter >= 965 AND x_counter <= 970) OR (x_counter >= 977 AND x_counter <= 982) OR (x_counter >= 986 AND x_counter <= 991) OR (x_counter >= 995 AND x_counter <= 1000) OR (x_counter >= 1004 AND x_counter <= 1018) OR (x_counter >= 1022 AND x_counter <= 1036) OR (x_counter >= 1040 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1063) OR (x_counter >= 1488 AND x_counter <= 1493) OR (x_counter >= 1500 AND x_counter <= 1505) OR (x_counter >= 1509 AND x_counter <= 1514) OR (x_counter >= 1518 AND x_counter <= 1523) OR (x_counter >= 1527 AND x_counter <= 1532) OR (x_counter >= 1542 AND x_counter <= 1556) OR (x_counter >= 1560 AND x_counter <= 1574) OR (x_counter >= 1578 AND x_counter <= 1592) OR (x_counter >= 1605 AND x_counter <= 1610) OR (x_counter >= 1617 AND x_counter <= 1622) OR (x_counter >= 1626 AND x_counter <= 1631) OR (x_counter >= 1635 AND x_counter <= 1640) OR (x_counter >= 1644 AND x_counter <= 1658) OR (x_counter >= 1662 AND x_counter <= 1676) OR (x_counter >= 1680 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1703)))
											OR	(y_counter = 391 AND ((x_counter >= 208 AND x_counter <= 213) OR (x_counter >= 220 AND x_counter <= 225) OR (x_counter >= 229 AND x_counter <= 234) OR (x_counter >= 238 AND x_counter <= 243) OR (x_counter >= 247 AND x_counter <= 252) OR (x_counter >= 262 AND x_counter <= 276) OR (x_counter >= 280 AND x_counter <= 294) OR (x_counter >= 298 AND x_counter <= 312) OR (x_counter >= 325 AND x_counter <= 330) OR (x_counter >= 337 AND x_counter <= 342) OR (x_counter >= 346 AND x_counter <= 351) OR (x_counter >= 355 AND x_counter <= 360) OR (x_counter >= 364 AND x_counter <= 378) OR (x_counter >= 382 AND x_counter <= 396) OR (x_counter >= 400 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 423) OR (x_counter >= 848 AND x_counter <= 853) OR (x_counter >= 860 AND x_counter <= 865) OR (x_counter >= 869 AND x_counter <= 874) OR (x_counter >= 878 AND x_counter <= 883) OR (x_counter >= 887 AND x_counter <= 892) OR (x_counter >= 902 AND x_counter <= 916) OR (x_counter >= 920 AND x_counter <= 934) OR (x_counter >= 938 AND x_counter <= 952) OR (x_counter >= 965 AND x_counter <= 970) OR (x_counter >= 977 AND x_counter <= 982) OR (x_counter >= 986 AND x_counter <= 991) OR (x_counter >= 995 AND x_counter <= 1000) OR (x_counter >= 1004 AND x_counter <= 1018) OR (x_counter >= 1022 AND x_counter <= 1036) OR (x_counter >= 1040 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1063) OR (x_counter >= 1488 AND x_counter <= 1493) OR (x_counter >= 1500 AND x_counter <= 1505) OR (x_counter >= 1509 AND x_counter <= 1514) OR (x_counter >= 1518 AND x_counter <= 1523) OR (x_counter >= 1527 AND x_counter <= 1532) OR (x_counter >= 1542 AND x_counter <= 1556) OR (x_counter >= 1560 AND x_counter <= 1574) OR (x_counter >= 1578 AND x_counter <= 1592) OR (x_counter >= 1605 AND x_counter <= 1610) OR (x_counter >= 1617 AND x_counter <= 1622) OR (x_counter >= 1626 AND x_counter <= 1631) OR (x_counter >= 1635 AND x_counter <= 1640) OR (x_counter >= 1644 AND x_counter <= 1658) OR (x_counter >= 1662 AND x_counter <= 1676) OR (x_counter >= 1680 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1703)))
											OR	(y_counter = 392 AND ((x_counter >= 364 AND x_counter <= 369) OR (x_counter >= 1004 AND x_counter <= 1009) OR (x_counter >= 1644 AND x_counter <= 1649)))
											OR	(y_counter = 393 AND ((x_counter >= 364 AND x_counter <= 369) OR (x_counter >= 1004 AND x_counter <= 1009) OR (x_counter >= 1644 AND x_counter <= 1649)))
											OR	(y_counter = 394 AND ((x_counter >= 364 AND x_counter <= 369) OR (x_counter >= 1004 AND x_counter <= 1009) OR (x_counter >= 1644 AND x_counter <= 1649)))
											OR	(y_counter = 395 AND ((x_counter >= 364 AND x_counter <= 369) OR (x_counter >= 1004 AND x_counter <= 1009) OR (x_counter >= 1644 AND x_counter <= 1649)))
											OR	(y_counter = 396 AND ((x_counter >= 364 AND x_counter <= 369) OR (x_counter >= 1004 AND x_counter <= 1009) OR (x_counter >= 1644 AND x_counter <= 1649)))
											OR	(y_counter = 397 AND ((x_counter >= 364 AND x_counter <= 369) OR (x_counter >= 1004 AND x_counter <= 1009) OR (x_counter >= 1644 AND x_counter <= 1649)))
											OR	(y_counter = 398 AND ((x_counter >= 364 AND x_counter <= 369) OR (x_counter >= 1004 AND x_counter <= 1009) OR (x_counter >= 1644 AND x_counter <= 1649)))
											OR	(y_counter = 399 AND ((x_counter >= 364 AND x_counter <= 369) OR (x_counter >= 1004 AND x_counter <= 1009) OR (x_counter >= 1644 AND x_counter <= 1649)))
											OR	(y_counter = 400 AND ((x_counter >= 364 AND x_counter <= 369) OR (x_counter >= 1004 AND x_counter <= 1009) OR (x_counter >= 1644 AND x_counter <= 1649)))
											OR	(y_counter = 402 AND ((x_counter >= 304 AND x_counter <= 309) OR (x_counter >= 313 AND x_counter <= 318) OR (x_counter >= 944 AND x_counter <= 949) OR (x_counter >= 953 AND x_counter <= 958) OR (x_counter >= 1584 AND x_counter <= 1589) OR (x_counter >= 1593 AND x_counter <= 1598)))
											OR	(y_counter = 403 AND ((x_counter >= 304 AND x_counter <= 309) OR (x_counter >= 313 AND x_counter <= 318) OR (x_counter >= 944 AND x_counter <= 949) OR (x_counter >= 953 AND x_counter <= 958) OR (x_counter >= 1584 AND x_counter <= 1589) OR (x_counter >= 1593 AND x_counter <= 1598)))
											OR	(y_counter = 404 AND ((x_counter >= 304 AND x_counter <= 309) OR (x_counter >= 313 AND x_counter <= 318) OR (x_counter >= 944 AND x_counter <= 949) OR (x_counter >= 953 AND x_counter <= 958) OR (x_counter >= 1584 AND x_counter <= 1589) OR (x_counter >= 1593 AND x_counter <= 1598)))
											OR	(y_counter = 405 AND ((x_counter >= 304 AND x_counter <= 309) OR (x_counter >= 313 AND x_counter <= 318) OR (x_counter >= 944 AND x_counter <= 949) OR (x_counter >= 953 AND x_counter <= 958) OR (x_counter >= 1584 AND x_counter <= 1589) OR (x_counter >= 1593 AND x_counter <= 1598)))
											OR	(y_counter = 406 AND ((x_counter >= 304 AND x_counter <= 309) OR (x_counter >= 313 AND x_counter <= 318) OR (x_counter >= 944 AND x_counter <= 949) OR (x_counter >= 953 AND x_counter <= 958) OR (x_counter >= 1584 AND x_counter <= 1589) OR (x_counter >= 1593 AND x_counter <= 1598)))
											OR	(y_counter = 407 AND ((x_counter >= 304 AND x_counter <= 309) OR (x_counter >= 313 AND x_counter <= 318) OR (x_counter >= 944 AND x_counter <= 949) OR (x_counter >= 953 AND x_counter <= 958) OR (x_counter >= 1584 AND x_counter <= 1589) OR (x_counter >= 1593 AND x_counter <= 1598)))
											OR	(y_counter = 408 AND ((x_counter >= 304 AND x_counter <= 309) OR (x_counter >= 944 AND x_counter <= 949) OR (x_counter >= 1584 AND x_counter <= 1589)))
											OR	(y_counter = 409 AND ((x_counter >= 304 AND x_counter <= 309) OR (x_counter >= 944 AND x_counter <= 949) OR (x_counter >= 1584 AND x_counter <= 1589)))
											OR	(y_counter = 410 AND ((x_counter >= 304 AND x_counter <= 309) OR (x_counter >= 944 AND x_counter <= 949) OR (x_counter >= 1584 AND x_counter <= 1589)))
											OR	(y_counter = 411 AND ((x_counter >= 196 AND x_counter <= 201) OR (x_counter >= 205 AND x_counter <= 210) OR (x_counter >= 214 AND x_counter <= 219) OR (x_counter >= 223 AND x_counter <= 228) OR (x_counter >= 232 AND x_counter <= 237) OR (x_counter >= 241 AND x_counter <= 246) OR (x_counter >= 250 AND x_counter <= 255) OR (x_counter >= 259 AND x_counter <= 264) OR (x_counter >= 268 AND x_counter <= 273) OR (x_counter >= 286 AND x_counter <= 300) OR (x_counter >= 304 AND x_counter <= 309) OR (x_counter >= 313 AND x_counter <= 318) OR (x_counter >= 322 AND x_counter <= 336) OR (x_counter >= 340 AND x_counter <= 354) OR (x_counter >= 358 AND x_counter <= 363) OR (x_counter >= 367 AND x_counter <= 372) OR (x_counter >= 376 AND x_counter <= 387) OR (x_counter >= 400 AND x_counter <= 423) OR (x_counter >= 427 AND x_counter <= 441) OR (x_counter >= 836 AND x_counter <= 841) OR (x_counter >= 845 AND x_counter <= 850) OR (x_counter >= 854 AND x_counter <= 859) OR (x_counter >= 863 AND x_counter <= 868) OR (x_counter >= 872 AND x_counter <= 877) OR (x_counter >= 881 AND x_counter <= 886) OR (x_counter >= 890 AND x_counter <= 895) OR (x_counter >= 899 AND x_counter <= 904) OR (x_counter >= 908 AND x_counter <= 913) OR (x_counter >= 926 AND x_counter <= 940) OR (x_counter >= 944 AND x_counter <= 949) OR (x_counter >= 953 AND x_counter <= 958) OR (x_counter >= 962 AND x_counter <= 976) OR (x_counter >= 980 AND x_counter <= 994) OR (x_counter >= 998 AND x_counter <= 1003) OR (x_counter >= 1007 AND x_counter <= 1012) OR (x_counter >= 1016 AND x_counter <= 1027) OR (x_counter >= 1040 AND x_counter <= 1063) OR (x_counter >= 1067 AND x_counter <= 1081) OR (x_counter >= 1476 AND x_counter <= 1481) OR (x_counter >= 1485 AND x_counter <= 1490) OR (x_counter >= 1494 AND x_counter <= 1499) OR (x_counter >= 1503 AND x_counter <= 1508) OR (x_counter >= 1512 AND x_counter <= 1517) OR (x_counter >= 1521 AND x_counter <= 1526) OR (x_counter >= 1530 AND x_counter <= 1535) OR (x_counter >= 1539 AND x_counter <= 1544) OR (x_counter >= 1548 AND x_counter <= 1553) OR (x_counter >= 1566 AND x_counter <= 1580) OR (x_counter >= 1584 AND x_counter <= 1589) OR (x_counter >= 1593 AND x_counter <= 1598) OR (x_counter >= 1602 AND x_counter <= 1616) OR (x_counter >= 1620 AND x_counter <= 1634) OR (x_counter >= 1638 AND x_counter <= 1643) OR (x_counter >= 1647 AND x_counter <= 1652) OR (x_counter >= 1656 AND x_counter <= 1667) OR (x_counter >= 1680 AND x_counter <= 1703) OR (x_counter >= 1707 AND x_counter <= 1721)))
											OR	(y_counter = 412 AND ((x_counter >= 196 AND x_counter <= 201) OR (x_counter >= 205 AND x_counter <= 210) OR (x_counter >= 214 AND x_counter <= 219) OR (x_counter >= 223 AND x_counter <= 228) OR (x_counter >= 232 AND x_counter <= 237) OR (x_counter >= 241 AND x_counter <= 246) OR (x_counter >= 250 AND x_counter <= 255) OR (x_counter >= 259 AND x_counter <= 264) OR (x_counter >= 268 AND x_counter <= 273) OR (x_counter >= 286 AND x_counter <= 300) OR (x_counter >= 304 AND x_counter <= 309) OR (x_counter >= 313 AND x_counter <= 318) OR (x_counter >= 322 AND x_counter <= 336) OR (x_counter >= 340 AND x_counter <= 354) OR (x_counter >= 358 AND x_counter <= 363) OR (x_counter >= 367 AND x_counter <= 372) OR (x_counter >= 376 AND x_counter <= 387) OR (x_counter >= 400 AND x_counter <= 423) OR (x_counter >= 427 AND x_counter <= 441) OR (x_counter >= 836 AND x_counter <= 841) OR (x_counter >= 845 AND x_counter <= 850) OR (x_counter >= 854 AND x_counter <= 859) OR (x_counter >= 863 AND x_counter <= 868) OR (x_counter >= 872 AND x_counter <= 877) OR (x_counter >= 881 AND x_counter <= 886) OR (x_counter >= 890 AND x_counter <= 895) OR (x_counter >= 899 AND x_counter <= 904) OR (x_counter >= 908 AND x_counter <= 913) OR (x_counter >= 926 AND x_counter <= 940) OR (x_counter >= 944 AND x_counter <= 949) OR (x_counter >= 953 AND x_counter <= 958) OR (x_counter >= 962 AND x_counter <= 976) OR (x_counter >= 980 AND x_counter <= 994) OR (x_counter >= 998 AND x_counter <= 1003) OR (x_counter >= 1007 AND x_counter <= 1012) OR (x_counter >= 1016 AND x_counter <= 1027) OR (x_counter >= 1040 AND x_counter <= 1063) OR (x_counter >= 1067 AND x_counter <= 1081) OR (x_counter >= 1476 AND x_counter <= 1481) OR (x_counter >= 1485 AND x_counter <= 1490) OR (x_counter >= 1494 AND x_counter <= 1499) OR (x_counter >= 1503 AND x_counter <= 1508) OR (x_counter >= 1512 AND x_counter <= 1517) OR (x_counter >= 1521 AND x_counter <= 1526) OR (x_counter >= 1530 AND x_counter <= 1535) OR (x_counter >= 1539 AND x_counter <= 1544) OR (x_counter >= 1548 AND x_counter <= 1553) OR (x_counter >= 1566 AND x_counter <= 1580) OR (x_counter >= 1584 AND x_counter <= 1589) OR (x_counter >= 1593 AND x_counter <= 1598) OR (x_counter >= 1602 AND x_counter <= 1616) OR (x_counter >= 1620 AND x_counter <= 1634) OR (x_counter >= 1638 AND x_counter <= 1643) OR (x_counter >= 1647 AND x_counter <= 1652) OR (x_counter >= 1656 AND x_counter <= 1667) OR (x_counter >= 1680 AND x_counter <= 1703) OR (x_counter >= 1707 AND x_counter <= 1721)))
											OR	(y_counter = 413 AND ((x_counter >= 196 AND x_counter <= 201) OR (x_counter >= 205 AND x_counter <= 210) OR (x_counter >= 214 AND x_counter <= 219) OR (x_counter >= 223 AND x_counter <= 228) OR (x_counter >= 232 AND x_counter <= 237) OR (x_counter >= 241 AND x_counter <= 246) OR (x_counter >= 250 AND x_counter <= 255) OR (x_counter >= 259 AND x_counter <= 264) OR (x_counter >= 268 AND x_counter <= 273) OR (x_counter >= 286 AND x_counter <= 300) OR (x_counter >= 304 AND x_counter <= 309) OR (x_counter >= 313 AND x_counter <= 318) OR (x_counter >= 322 AND x_counter <= 336) OR (x_counter >= 340 AND x_counter <= 354) OR (x_counter >= 358 AND x_counter <= 363) OR (x_counter >= 367 AND x_counter <= 372) OR (x_counter >= 376 AND x_counter <= 387) OR (x_counter >= 400 AND x_counter <= 423) OR (x_counter >= 427 AND x_counter <= 441) OR (x_counter >= 836 AND x_counter <= 841) OR (x_counter >= 845 AND x_counter <= 850) OR (x_counter >= 854 AND x_counter <= 859) OR (x_counter >= 863 AND x_counter <= 868) OR (x_counter >= 872 AND x_counter <= 877) OR (x_counter >= 881 AND x_counter <= 886) OR (x_counter >= 890 AND x_counter <= 895) OR (x_counter >= 899 AND x_counter <= 904) OR (x_counter >= 908 AND x_counter <= 913) OR (x_counter >= 926 AND x_counter <= 940) OR (x_counter >= 944 AND x_counter <= 949) OR (x_counter >= 953 AND x_counter <= 958) OR (x_counter >= 962 AND x_counter <= 976) OR (x_counter >= 980 AND x_counter <= 994) OR (x_counter >= 998 AND x_counter <= 1003) OR (x_counter >= 1007 AND x_counter <= 1012) OR (x_counter >= 1016 AND x_counter <= 1027) OR (x_counter >= 1040 AND x_counter <= 1063) OR (x_counter >= 1067 AND x_counter <= 1081) OR (x_counter >= 1476 AND x_counter <= 1481) OR (x_counter >= 1485 AND x_counter <= 1490) OR (x_counter >= 1494 AND x_counter <= 1499) OR (x_counter >= 1503 AND x_counter <= 1508) OR (x_counter >= 1512 AND x_counter <= 1517) OR (x_counter >= 1521 AND x_counter <= 1526) OR (x_counter >= 1530 AND x_counter <= 1535) OR (x_counter >= 1539 AND x_counter <= 1544) OR (x_counter >= 1548 AND x_counter <= 1553) OR (x_counter >= 1566 AND x_counter <= 1580) OR (x_counter >= 1584 AND x_counter <= 1589) OR (x_counter >= 1593 AND x_counter <= 1598) OR (x_counter >= 1602 AND x_counter <= 1616) OR (x_counter >= 1620 AND x_counter <= 1634) OR (x_counter >= 1638 AND x_counter <= 1643) OR (x_counter >= 1647 AND x_counter <= 1652) OR (x_counter >= 1656 AND x_counter <= 1667) OR (x_counter >= 1680 AND x_counter <= 1703) OR (x_counter >= 1707 AND x_counter <= 1721)))
											OR	(y_counter = 414 AND ((x_counter >= 196 AND x_counter <= 201) OR (x_counter >= 205 AND x_counter <= 210) OR (x_counter >= 214 AND x_counter <= 219) OR (x_counter >= 223 AND x_counter <= 228) OR (x_counter >= 232 AND x_counter <= 237) OR (x_counter >= 241 AND x_counter <= 246) OR (x_counter >= 250 AND x_counter <= 255) OR (x_counter >= 259 AND x_counter <= 264) OR (x_counter >= 268 AND x_counter <= 273) OR (x_counter >= 286 AND x_counter <= 300) OR (x_counter >= 304 AND x_counter <= 309) OR (x_counter >= 313 AND x_counter <= 318) OR (x_counter >= 322 AND x_counter <= 336) OR (x_counter >= 340 AND x_counter <= 354) OR (x_counter >= 358 AND x_counter <= 363) OR (x_counter >= 367 AND x_counter <= 372) OR (x_counter >= 376 AND x_counter <= 387) OR (x_counter >= 400 AND x_counter <= 423) OR (x_counter >= 427 AND x_counter <= 441) OR (x_counter >= 836 AND x_counter <= 841) OR (x_counter >= 845 AND x_counter <= 850) OR (x_counter >= 854 AND x_counter <= 859) OR (x_counter >= 863 AND x_counter <= 868) OR (x_counter >= 872 AND x_counter <= 877) OR (x_counter >= 881 AND x_counter <= 886) OR (x_counter >= 890 AND x_counter <= 895) OR (x_counter >= 899 AND x_counter <= 904) OR (x_counter >= 908 AND x_counter <= 913) OR (x_counter >= 926 AND x_counter <= 940) OR (x_counter >= 944 AND x_counter <= 949) OR (x_counter >= 953 AND x_counter <= 958) OR (x_counter >= 962 AND x_counter <= 976) OR (x_counter >= 980 AND x_counter <= 994) OR (x_counter >= 998 AND x_counter <= 1003) OR (x_counter >= 1007 AND x_counter <= 1012) OR (x_counter >= 1016 AND x_counter <= 1027) OR (x_counter >= 1040 AND x_counter <= 1063) OR (x_counter >= 1067 AND x_counter <= 1081) OR (x_counter >= 1476 AND x_counter <= 1481) OR (x_counter >= 1485 AND x_counter <= 1490) OR (x_counter >= 1494 AND x_counter <= 1499) OR (x_counter >= 1503 AND x_counter <= 1508) OR (x_counter >= 1512 AND x_counter <= 1517) OR (x_counter >= 1521 AND x_counter <= 1526) OR (x_counter >= 1530 AND x_counter <= 1535) OR (x_counter >= 1539 AND x_counter <= 1544) OR (x_counter >= 1548 AND x_counter <= 1553) OR (x_counter >= 1566 AND x_counter <= 1580) OR (x_counter >= 1584 AND x_counter <= 1589) OR (x_counter >= 1593 AND x_counter <= 1598) OR (x_counter >= 1602 AND x_counter <= 1616) OR (x_counter >= 1620 AND x_counter <= 1634) OR (x_counter >= 1638 AND x_counter <= 1643) OR (x_counter >= 1647 AND x_counter <= 1652) OR (x_counter >= 1656 AND x_counter <= 1667) OR (x_counter >= 1680 AND x_counter <= 1703) OR (x_counter >= 1707 AND x_counter <= 1721)))
											OR	(y_counter = 415 AND ((x_counter >= 196 AND x_counter <= 201) OR (x_counter >= 205 AND x_counter <= 210) OR (x_counter >= 214 AND x_counter <= 219) OR (x_counter >= 223 AND x_counter <= 228) OR (x_counter >= 232 AND x_counter <= 237) OR (x_counter >= 241 AND x_counter <= 246) OR (x_counter >= 250 AND x_counter <= 255) OR (x_counter >= 259 AND x_counter <= 264) OR (x_counter >= 268 AND x_counter <= 273) OR (x_counter >= 286 AND x_counter <= 300) OR (x_counter >= 304 AND x_counter <= 309) OR (x_counter >= 313 AND x_counter <= 318) OR (x_counter >= 322 AND x_counter <= 336) OR (x_counter >= 340 AND x_counter <= 354) OR (x_counter >= 358 AND x_counter <= 363) OR (x_counter >= 367 AND x_counter <= 372) OR (x_counter >= 376 AND x_counter <= 387) OR (x_counter >= 400 AND x_counter <= 423) OR (x_counter >= 427 AND x_counter <= 441) OR (x_counter >= 836 AND x_counter <= 841) OR (x_counter >= 845 AND x_counter <= 850) OR (x_counter >= 854 AND x_counter <= 859) OR (x_counter >= 863 AND x_counter <= 868) OR (x_counter >= 872 AND x_counter <= 877) OR (x_counter >= 881 AND x_counter <= 886) OR (x_counter >= 890 AND x_counter <= 895) OR (x_counter >= 899 AND x_counter <= 904) OR (x_counter >= 908 AND x_counter <= 913) OR (x_counter >= 926 AND x_counter <= 940) OR (x_counter >= 944 AND x_counter <= 949) OR (x_counter >= 953 AND x_counter <= 958) OR (x_counter >= 962 AND x_counter <= 976) OR (x_counter >= 980 AND x_counter <= 994) OR (x_counter >= 998 AND x_counter <= 1003) OR (x_counter >= 1007 AND x_counter <= 1012) OR (x_counter >= 1016 AND x_counter <= 1027) OR (x_counter >= 1040 AND x_counter <= 1063) OR (x_counter >= 1067 AND x_counter <= 1081) OR (x_counter >= 1476 AND x_counter <= 1481) OR (x_counter >= 1485 AND x_counter <= 1490) OR (x_counter >= 1494 AND x_counter <= 1499) OR (x_counter >= 1503 AND x_counter <= 1508) OR (x_counter >= 1512 AND x_counter <= 1517) OR (x_counter >= 1521 AND x_counter <= 1526) OR (x_counter >= 1530 AND x_counter <= 1535) OR (x_counter >= 1539 AND x_counter <= 1544) OR (x_counter >= 1548 AND x_counter <= 1553) OR (x_counter >= 1566 AND x_counter <= 1580) OR (x_counter >= 1584 AND x_counter <= 1589) OR (x_counter >= 1593 AND x_counter <= 1598) OR (x_counter >= 1602 AND x_counter <= 1616) OR (x_counter >= 1620 AND x_counter <= 1634) OR (x_counter >= 1638 AND x_counter <= 1643) OR (x_counter >= 1647 AND x_counter <= 1652) OR (x_counter >= 1656 AND x_counter <= 1667) OR (x_counter >= 1680 AND x_counter <= 1703) OR (x_counter >= 1707 AND x_counter <= 1721)))
											OR	(y_counter = 416 AND ((x_counter >= 196 AND x_counter <= 201) OR (x_counter >= 205 AND x_counter <= 210) OR (x_counter >= 214 AND x_counter <= 219) OR (x_counter >= 223 AND x_counter <= 228) OR (x_counter >= 232 AND x_counter <= 237) OR (x_counter >= 241 AND x_counter <= 246) OR (x_counter >= 250 AND x_counter <= 255) OR (x_counter >= 259 AND x_counter <= 264) OR (x_counter >= 268 AND x_counter <= 273) OR (x_counter >= 286 AND x_counter <= 300) OR (x_counter >= 304 AND x_counter <= 309) OR (x_counter >= 313 AND x_counter <= 318) OR (x_counter >= 322 AND x_counter <= 336) OR (x_counter >= 340 AND x_counter <= 354) OR (x_counter >= 358 AND x_counter <= 363) OR (x_counter >= 367 AND x_counter <= 372) OR (x_counter >= 376 AND x_counter <= 387) OR (x_counter >= 400 AND x_counter <= 423) OR (x_counter >= 427 AND x_counter <= 441) OR (x_counter >= 836 AND x_counter <= 841) OR (x_counter >= 845 AND x_counter <= 850) OR (x_counter >= 854 AND x_counter <= 859) OR (x_counter >= 863 AND x_counter <= 868) OR (x_counter >= 872 AND x_counter <= 877) OR (x_counter >= 881 AND x_counter <= 886) OR (x_counter >= 890 AND x_counter <= 895) OR (x_counter >= 899 AND x_counter <= 904) OR (x_counter >= 908 AND x_counter <= 913) OR (x_counter >= 926 AND x_counter <= 940) OR (x_counter >= 944 AND x_counter <= 949) OR (x_counter >= 953 AND x_counter <= 958) OR (x_counter >= 962 AND x_counter <= 976) OR (x_counter >= 980 AND x_counter <= 994) OR (x_counter >= 998 AND x_counter <= 1003) OR (x_counter >= 1007 AND x_counter <= 1012) OR (x_counter >= 1016 AND x_counter <= 1027) OR (x_counter >= 1040 AND x_counter <= 1063) OR (x_counter >= 1067 AND x_counter <= 1081) OR (x_counter >= 1476 AND x_counter <= 1481) OR (x_counter >= 1485 AND x_counter <= 1490) OR (x_counter >= 1494 AND x_counter <= 1499) OR (x_counter >= 1503 AND x_counter <= 1508) OR (x_counter >= 1512 AND x_counter <= 1517) OR (x_counter >= 1521 AND x_counter <= 1526) OR (x_counter >= 1530 AND x_counter <= 1535) OR (x_counter >= 1539 AND x_counter <= 1544) OR (x_counter >= 1548 AND x_counter <= 1553) OR (x_counter >= 1566 AND x_counter <= 1580) OR (x_counter >= 1584 AND x_counter <= 1589) OR (x_counter >= 1593 AND x_counter <= 1598) OR (x_counter >= 1602 AND x_counter <= 1616) OR (x_counter >= 1620 AND x_counter <= 1634) OR (x_counter >= 1638 AND x_counter <= 1643) OR (x_counter >= 1647 AND x_counter <= 1652) OR (x_counter >= 1656 AND x_counter <= 1667) OR (x_counter >= 1680 AND x_counter <= 1703) OR (x_counter >= 1707 AND x_counter <= 1721)))
											OR	(y_counter = 417 AND ((x_counter >= 196 AND x_counter <= 201) OR (x_counter >= 205 AND x_counter <= 210) OR (x_counter >= 214 AND x_counter <= 219) OR (x_counter >= 223 AND x_counter <= 228) OR (x_counter >= 232 AND x_counter <= 237) OR (x_counter >= 241 AND x_counter <= 246) OR (x_counter >= 250 AND x_counter <= 255) OR (x_counter >= 259 AND x_counter <= 264) OR (x_counter >= 268 AND x_counter <= 273) OR (x_counter >= 295 AND x_counter <= 300) OR (x_counter >= 304 AND x_counter <= 309) OR (x_counter >= 313 AND x_counter <= 318) OR (x_counter >= 322 AND x_counter <= 327) OR (x_counter >= 331 AND x_counter <= 336) OR (x_counter >= 340 AND x_counter <= 345) OR (x_counter >= 349 AND x_counter <= 354) OR (x_counter >= 358 AND x_counter <= 363) OR (x_counter >= 367 AND x_counter <= 372) OR (x_counter >= 376 AND x_counter <= 381) OR (x_counter >= 400 AND x_counter <= 405) OR (x_counter >= 409 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 423) OR (x_counter >= 427 AND x_counter <= 432) OR (x_counter >= 436 AND x_counter <= 441) OR (x_counter >= 836 AND x_counter <= 841) OR (x_counter >= 845 AND x_counter <= 850) OR (x_counter >= 854 AND x_counter <= 859) OR (x_counter >= 863 AND x_counter <= 868) OR (x_counter >= 872 AND x_counter <= 877) OR (x_counter >= 881 AND x_counter <= 886) OR (x_counter >= 890 AND x_counter <= 895) OR (x_counter >= 899 AND x_counter <= 904) OR (x_counter >= 908 AND x_counter <= 913) OR (x_counter >= 935 AND x_counter <= 940) OR (x_counter >= 944 AND x_counter <= 949) OR (x_counter >= 953 AND x_counter <= 958) OR (x_counter >= 962 AND x_counter <= 967) OR (x_counter >= 971 AND x_counter <= 976) OR (x_counter >= 980 AND x_counter <= 985) OR (x_counter >= 989 AND x_counter <= 994) OR (x_counter >= 998 AND x_counter <= 1003) OR (x_counter >= 1007 AND x_counter <= 1012) OR (x_counter >= 1016 AND x_counter <= 1021) OR (x_counter >= 1040 AND x_counter <= 1045) OR (x_counter >= 1049 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1063) OR (x_counter >= 1067 AND x_counter <= 1072) OR (x_counter >= 1076 AND x_counter <= 1081) OR (x_counter >= 1476 AND x_counter <= 1481) OR (x_counter >= 1485 AND x_counter <= 1490) OR (x_counter >= 1494 AND x_counter <= 1499) OR (x_counter >= 1503 AND x_counter <= 1508) OR (x_counter >= 1512 AND x_counter <= 1517) OR (x_counter >= 1521 AND x_counter <= 1526) OR (x_counter >= 1530 AND x_counter <= 1535) OR (x_counter >= 1539 AND x_counter <= 1544) OR (x_counter >= 1548 AND x_counter <= 1553) OR (x_counter >= 1575 AND x_counter <= 1580) OR (x_counter >= 1584 AND x_counter <= 1589) OR (x_counter >= 1593 AND x_counter <= 1598) OR (x_counter >= 1602 AND x_counter <= 1607) OR (x_counter >= 1611 AND x_counter <= 1616) OR (x_counter >= 1620 AND x_counter <= 1625) OR (x_counter >= 1629 AND x_counter <= 1634) OR (x_counter >= 1638 AND x_counter <= 1643) OR (x_counter >= 1647 AND x_counter <= 1652) OR (x_counter >= 1656 AND x_counter <= 1661) OR (x_counter >= 1680 AND x_counter <= 1685) OR (x_counter >= 1689 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1703) OR (x_counter >= 1707 AND x_counter <= 1712) OR (x_counter >= 1716 AND x_counter <= 1721)))
											OR	(y_counter = 418 AND ((x_counter >= 196 AND x_counter <= 201) OR (x_counter >= 205 AND x_counter <= 210) OR (x_counter >= 214 AND x_counter <= 219) OR (x_counter >= 223 AND x_counter <= 228) OR (x_counter >= 232 AND x_counter <= 237) OR (x_counter >= 241 AND x_counter <= 246) OR (x_counter >= 250 AND x_counter <= 255) OR (x_counter >= 259 AND x_counter <= 264) OR (x_counter >= 268 AND x_counter <= 273) OR (x_counter >= 295 AND x_counter <= 300) OR (x_counter >= 304 AND x_counter <= 309) OR (x_counter >= 313 AND x_counter <= 318) OR (x_counter >= 322 AND x_counter <= 327) OR (x_counter >= 331 AND x_counter <= 336) OR (x_counter >= 340 AND x_counter <= 345) OR (x_counter >= 349 AND x_counter <= 354) OR (x_counter >= 358 AND x_counter <= 363) OR (x_counter >= 367 AND x_counter <= 372) OR (x_counter >= 376 AND x_counter <= 381) OR (x_counter >= 400 AND x_counter <= 405) OR (x_counter >= 409 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 423) OR (x_counter >= 427 AND x_counter <= 432) OR (x_counter >= 436 AND x_counter <= 441) OR (x_counter >= 836 AND x_counter <= 841) OR (x_counter >= 845 AND x_counter <= 850) OR (x_counter >= 854 AND x_counter <= 859) OR (x_counter >= 863 AND x_counter <= 868) OR (x_counter >= 872 AND x_counter <= 877) OR (x_counter >= 881 AND x_counter <= 886) OR (x_counter >= 890 AND x_counter <= 895) OR (x_counter >= 899 AND x_counter <= 904) OR (x_counter >= 908 AND x_counter <= 913) OR (x_counter >= 935 AND x_counter <= 940) OR (x_counter >= 944 AND x_counter <= 949) OR (x_counter >= 953 AND x_counter <= 958) OR (x_counter >= 962 AND x_counter <= 967) OR (x_counter >= 971 AND x_counter <= 976) OR (x_counter >= 980 AND x_counter <= 985) OR (x_counter >= 989 AND x_counter <= 994) OR (x_counter >= 998 AND x_counter <= 1003) OR (x_counter >= 1007 AND x_counter <= 1012) OR (x_counter >= 1016 AND x_counter <= 1021) OR (x_counter >= 1040 AND x_counter <= 1045) OR (x_counter >= 1049 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1063) OR (x_counter >= 1067 AND x_counter <= 1072) OR (x_counter >= 1076 AND x_counter <= 1081) OR (x_counter >= 1476 AND x_counter <= 1481) OR (x_counter >= 1485 AND x_counter <= 1490) OR (x_counter >= 1494 AND x_counter <= 1499) OR (x_counter >= 1503 AND x_counter <= 1508) OR (x_counter >= 1512 AND x_counter <= 1517) OR (x_counter >= 1521 AND x_counter <= 1526) OR (x_counter >= 1530 AND x_counter <= 1535) OR (x_counter >= 1539 AND x_counter <= 1544) OR (x_counter >= 1548 AND x_counter <= 1553) OR (x_counter >= 1575 AND x_counter <= 1580) OR (x_counter >= 1584 AND x_counter <= 1589) OR (x_counter >= 1593 AND x_counter <= 1598) OR (x_counter >= 1602 AND x_counter <= 1607) OR (x_counter >= 1611 AND x_counter <= 1616) OR (x_counter >= 1620 AND x_counter <= 1625) OR (x_counter >= 1629 AND x_counter <= 1634) OR (x_counter >= 1638 AND x_counter <= 1643) OR (x_counter >= 1647 AND x_counter <= 1652) OR (x_counter >= 1656 AND x_counter <= 1661) OR (x_counter >= 1680 AND x_counter <= 1685) OR (x_counter >= 1689 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1703) OR (x_counter >= 1707 AND x_counter <= 1712) OR (x_counter >= 1716 AND x_counter <= 1721)))
											OR	(y_counter = 419 AND ((x_counter >= 196 AND x_counter <= 201) OR (x_counter >= 205 AND x_counter <= 210) OR (x_counter >= 214 AND x_counter <= 219) OR (x_counter >= 223 AND x_counter <= 228) OR (x_counter >= 232 AND x_counter <= 237) OR (x_counter >= 241 AND x_counter <= 246) OR (x_counter >= 250 AND x_counter <= 255) OR (x_counter >= 259 AND x_counter <= 264) OR (x_counter >= 268 AND x_counter <= 273) OR (x_counter >= 295 AND x_counter <= 300) OR (x_counter >= 304 AND x_counter <= 309) OR (x_counter >= 313 AND x_counter <= 318) OR (x_counter >= 322 AND x_counter <= 327) OR (x_counter >= 331 AND x_counter <= 336) OR (x_counter >= 340 AND x_counter <= 345) OR (x_counter >= 349 AND x_counter <= 354) OR (x_counter >= 358 AND x_counter <= 363) OR (x_counter >= 367 AND x_counter <= 372) OR (x_counter >= 376 AND x_counter <= 381) OR (x_counter >= 400 AND x_counter <= 405) OR (x_counter >= 409 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 423) OR (x_counter >= 427 AND x_counter <= 432) OR (x_counter >= 436 AND x_counter <= 441) OR (x_counter >= 836 AND x_counter <= 841) OR (x_counter >= 845 AND x_counter <= 850) OR (x_counter >= 854 AND x_counter <= 859) OR (x_counter >= 863 AND x_counter <= 868) OR (x_counter >= 872 AND x_counter <= 877) OR (x_counter >= 881 AND x_counter <= 886) OR (x_counter >= 890 AND x_counter <= 895) OR (x_counter >= 899 AND x_counter <= 904) OR (x_counter >= 908 AND x_counter <= 913) OR (x_counter >= 935 AND x_counter <= 940) OR (x_counter >= 944 AND x_counter <= 949) OR (x_counter >= 953 AND x_counter <= 958) OR (x_counter >= 962 AND x_counter <= 967) OR (x_counter >= 971 AND x_counter <= 976) OR (x_counter >= 980 AND x_counter <= 985) OR (x_counter >= 989 AND x_counter <= 994) OR (x_counter >= 998 AND x_counter <= 1003) OR (x_counter >= 1007 AND x_counter <= 1012) OR (x_counter >= 1016 AND x_counter <= 1021) OR (x_counter >= 1040 AND x_counter <= 1045) OR (x_counter >= 1049 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1063) OR (x_counter >= 1067 AND x_counter <= 1072) OR (x_counter >= 1076 AND x_counter <= 1081) OR (x_counter >= 1476 AND x_counter <= 1481) OR (x_counter >= 1485 AND x_counter <= 1490) OR (x_counter >= 1494 AND x_counter <= 1499) OR (x_counter >= 1503 AND x_counter <= 1508) OR (x_counter >= 1512 AND x_counter <= 1517) OR (x_counter >= 1521 AND x_counter <= 1526) OR (x_counter >= 1530 AND x_counter <= 1535) OR (x_counter >= 1539 AND x_counter <= 1544) OR (x_counter >= 1548 AND x_counter <= 1553) OR (x_counter >= 1575 AND x_counter <= 1580) OR (x_counter >= 1584 AND x_counter <= 1589) OR (x_counter >= 1593 AND x_counter <= 1598) OR (x_counter >= 1602 AND x_counter <= 1607) OR (x_counter >= 1611 AND x_counter <= 1616) OR (x_counter >= 1620 AND x_counter <= 1625) OR (x_counter >= 1629 AND x_counter <= 1634) OR (x_counter >= 1638 AND x_counter <= 1643) OR (x_counter >= 1647 AND x_counter <= 1652) OR (x_counter >= 1656 AND x_counter <= 1661) OR (x_counter >= 1680 AND x_counter <= 1685) OR (x_counter >= 1689 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1703) OR (x_counter >= 1707 AND x_counter <= 1712) OR (x_counter >= 1716 AND x_counter <= 1721)))
											OR	(y_counter = 420 AND ((x_counter >= 196 AND x_counter <= 201) OR (x_counter >= 205 AND x_counter <= 210) OR (x_counter >= 214 AND x_counter <= 219) OR (x_counter >= 223 AND x_counter <= 228) OR (x_counter >= 232 AND x_counter <= 237) OR (x_counter >= 241 AND x_counter <= 246) OR (x_counter >= 250 AND x_counter <= 255) OR (x_counter >= 259 AND x_counter <= 264) OR (x_counter >= 268 AND x_counter <= 273) OR (x_counter >= 286 AND x_counter <= 300) OR (x_counter >= 304 AND x_counter <= 309) OR (x_counter >= 313 AND x_counter <= 318) OR (x_counter >= 322 AND x_counter <= 327) OR (x_counter >= 331 AND x_counter <= 336) OR (x_counter >= 340 AND x_counter <= 345) OR (x_counter >= 349 AND x_counter <= 354) OR (x_counter >= 358 AND x_counter <= 363) OR (x_counter >= 367 AND x_counter <= 372) OR (x_counter >= 376 AND x_counter <= 381) OR (x_counter >= 400 AND x_counter <= 405) OR (x_counter >= 409 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 423) OR (x_counter >= 427 AND x_counter <= 441) OR (x_counter >= 836 AND x_counter <= 841) OR (x_counter >= 845 AND x_counter <= 850) OR (x_counter >= 854 AND x_counter <= 859) OR (x_counter >= 863 AND x_counter <= 868) OR (x_counter >= 872 AND x_counter <= 877) OR (x_counter >= 881 AND x_counter <= 886) OR (x_counter >= 890 AND x_counter <= 895) OR (x_counter >= 899 AND x_counter <= 904) OR (x_counter >= 908 AND x_counter <= 913) OR (x_counter >= 926 AND x_counter <= 940) OR (x_counter >= 944 AND x_counter <= 949) OR (x_counter >= 953 AND x_counter <= 958) OR (x_counter >= 962 AND x_counter <= 967) OR (x_counter >= 971 AND x_counter <= 976) OR (x_counter >= 980 AND x_counter <= 985) OR (x_counter >= 989 AND x_counter <= 994) OR (x_counter >= 998 AND x_counter <= 1003) OR (x_counter >= 1007 AND x_counter <= 1012) OR (x_counter >= 1016 AND x_counter <= 1021) OR (x_counter >= 1040 AND x_counter <= 1045) OR (x_counter >= 1049 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1063) OR (x_counter >= 1067 AND x_counter <= 1081) OR (x_counter >= 1476 AND x_counter <= 1481) OR (x_counter >= 1485 AND x_counter <= 1490) OR (x_counter >= 1494 AND x_counter <= 1499) OR (x_counter >= 1503 AND x_counter <= 1508) OR (x_counter >= 1512 AND x_counter <= 1517) OR (x_counter >= 1521 AND x_counter <= 1526) OR (x_counter >= 1530 AND x_counter <= 1535) OR (x_counter >= 1539 AND x_counter <= 1544) OR (x_counter >= 1548 AND x_counter <= 1553) OR (x_counter >= 1566 AND x_counter <= 1580) OR (x_counter >= 1584 AND x_counter <= 1589) OR (x_counter >= 1593 AND x_counter <= 1598) OR (x_counter >= 1602 AND x_counter <= 1607) OR (x_counter >= 1611 AND x_counter <= 1616) OR (x_counter >= 1620 AND x_counter <= 1625) OR (x_counter >= 1629 AND x_counter <= 1634) OR (x_counter >= 1638 AND x_counter <= 1643) OR (x_counter >= 1647 AND x_counter <= 1652) OR (x_counter >= 1656 AND x_counter <= 1661) OR (x_counter >= 1680 AND x_counter <= 1685) OR (x_counter >= 1689 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1703) OR (x_counter >= 1707 AND x_counter <= 1721)))
											OR	(y_counter = 421 AND ((x_counter >= 196 AND x_counter <= 201) OR (x_counter >= 205 AND x_counter <= 210) OR (x_counter >= 214 AND x_counter <= 219) OR (x_counter >= 223 AND x_counter <= 228) OR (x_counter >= 232 AND x_counter <= 237) OR (x_counter >= 241 AND x_counter <= 246) OR (x_counter >= 250 AND x_counter <= 255) OR (x_counter >= 259 AND x_counter <= 264) OR (x_counter >= 268 AND x_counter <= 273) OR (x_counter >= 286 AND x_counter <= 300) OR (x_counter >= 304 AND x_counter <= 309) OR (x_counter >= 313 AND x_counter <= 318) OR (x_counter >= 322 AND x_counter <= 327) OR (x_counter >= 331 AND x_counter <= 336) OR (x_counter >= 340 AND x_counter <= 345) OR (x_counter >= 349 AND x_counter <= 354) OR (x_counter >= 358 AND x_counter <= 363) OR (x_counter >= 367 AND x_counter <= 372) OR (x_counter >= 376 AND x_counter <= 381) OR (x_counter >= 400 AND x_counter <= 405) OR (x_counter >= 409 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 423) OR (x_counter >= 427 AND x_counter <= 441) OR (x_counter >= 836 AND x_counter <= 841) OR (x_counter >= 845 AND x_counter <= 850) OR (x_counter >= 854 AND x_counter <= 859) OR (x_counter >= 863 AND x_counter <= 868) OR (x_counter >= 872 AND x_counter <= 877) OR (x_counter >= 881 AND x_counter <= 886) OR (x_counter >= 890 AND x_counter <= 895) OR (x_counter >= 899 AND x_counter <= 904) OR (x_counter >= 908 AND x_counter <= 913) OR (x_counter >= 926 AND x_counter <= 940) OR (x_counter >= 944 AND x_counter <= 949) OR (x_counter >= 953 AND x_counter <= 958) OR (x_counter >= 962 AND x_counter <= 967) OR (x_counter >= 971 AND x_counter <= 976) OR (x_counter >= 980 AND x_counter <= 985) OR (x_counter >= 989 AND x_counter <= 994) OR (x_counter >= 998 AND x_counter <= 1003) OR (x_counter >= 1007 AND x_counter <= 1012) OR (x_counter >= 1016 AND x_counter <= 1021) OR (x_counter >= 1040 AND x_counter <= 1045) OR (x_counter >= 1049 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1063) OR (x_counter >= 1067 AND x_counter <= 1081) OR (x_counter >= 1476 AND x_counter <= 1481) OR (x_counter >= 1485 AND x_counter <= 1490) OR (x_counter >= 1494 AND x_counter <= 1499) OR (x_counter >= 1503 AND x_counter <= 1508) OR (x_counter >= 1512 AND x_counter <= 1517) OR (x_counter >= 1521 AND x_counter <= 1526) OR (x_counter >= 1530 AND x_counter <= 1535) OR (x_counter >= 1539 AND x_counter <= 1544) OR (x_counter >= 1548 AND x_counter <= 1553) OR (x_counter >= 1566 AND x_counter <= 1580) OR (x_counter >= 1584 AND x_counter <= 1589) OR (x_counter >= 1593 AND x_counter <= 1598) OR (x_counter >= 1602 AND x_counter <= 1607) OR (x_counter >= 1611 AND x_counter <= 1616) OR (x_counter >= 1620 AND x_counter <= 1625) OR (x_counter >= 1629 AND x_counter <= 1634) OR (x_counter >= 1638 AND x_counter <= 1643) OR (x_counter >= 1647 AND x_counter <= 1652) OR (x_counter >= 1656 AND x_counter <= 1661) OR (x_counter >= 1680 AND x_counter <= 1685) OR (x_counter >= 1689 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1703) OR (x_counter >= 1707 AND x_counter <= 1721)))
											OR	(y_counter = 422 AND ((x_counter >= 196 AND x_counter <= 201) OR (x_counter >= 205 AND x_counter <= 210) OR (x_counter >= 214 AND x_counter <= 219) OR (x_counter >= 223 AND x_counter <= 228) OR (x_counter >= 232 AND x_counter <= 237) OR (x_counter >= 241 AND x_counter <= 246) OR (x_counter >= 250 AND x_counter <= 255) OR (x_counter >= 259 AND x_counter <= 264) OR (x_counter >= 268 AND x_counter <= 273) OR (x_counter >= 286 AND x_counter <= 300) OR (x_counter >= 304 AND x_counter <= 309) OR (x_counter >= 313 AND x_counter <= 318) OR (x_counter >= 322 AND x_counter <= 327) OR (x_counter >= 331 AND x_counter <= 336) OR (x_counter >= 340 AND x_counter <= 345) OR (x_counter >= 349 AND x_counter <= 354) OR (x_counter >= 358 AND x_counter <= 363) OR (x_counter >= 367 AND x_counter <= 372) OR (x_counter >= 376 AND x_counter <= 381) OR (x_counter >= 400 AND x_counter <= 405) OR (x_counter >= 409 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 423) OR (x_counter >= 427 AND x_counter <= 441) OR (x_counter >= 836 AND x_counter <= 841) OR (x_counter >= 845 AND x_counter <= 850) OR (x_counter >= 854 AND x_counter <= 859) OR (x_counter >= 863 AND x_counter <= 868) OR (x_counter >= 872 AND x_counter <= 877) OR (x_counter >= 881 AND x_counter <= 886) OR (x_counter >= 890 AND x_counter <= 895) OR (x_counter >= 899 AND x_counter <= 904) OR (x_counter >= 908 AND x_counter <= 913) OR (x_counter >= 926 AND x_counter <= 940) OR (x_counter >= 944 AND x_counter <= 949) OR (x_counter >= 953 AND x_counter <= 958) OR (x_counter >= 962 AND x_counter <= 967) OR (x_counter >= 971 AND x_counter <= 976) OR (x_counter >= 980 AND x_counter <= 985) OR (x_counter >= 989 AND x_counter <= 994) OR (x_counter >= 998 AND x_counter <= 1003) OR (x_counter >= 1007 AND x_counter <= 1012) OR (x_counter >= 1016 AND x_counter <= 1021) OR (x_counter >= 1040 AND x_counter <= 1045) OR (x_counter >= 1049 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1063) OR (x_counter >= 1067 AND x_counter <= 1081) OR (x_counter >= 1476 AND x_counter <= 1481) OR (x_counter >= 1485 AND x_counter <= 1490) OR (x_counter >= 1494 AND x_counter <= 1499) OR (x_counter >= 1503 AND x_counter <= 1508) OR (x_counter >= 1512 AND x_counter <= 1517) OR (x_counter >= 1521 AND x_counter <= 1526) OR (x_counter >= 1530 AND x_counter <= 1535) OR (x_counter >= 1539 AND x_counter <= 1544) OR (x_counter >= 1548 AND x_counter <= 1553) OR (x_counter >= 1566 AND x_counter <= 1580) OR (x_counter >= 1584 AND x_counter <= 1589) OR (x_counter >= 1593 AND x_counter <= 1598) OR (x_counter >= 1602 AND x_counter <= 1607) OR (x_counter >= 1611 AND x_counter <= 1616) OR (x_counter >= 1620 AND x_counter <= 1625) OR (x_counter >= 1629 AND x_counter <= 1634) OR (x_counter >= 1638 AND x_counter <= 1643) OR (x_counter >= 1647 AND x_counter <= 1652) OR (x_counter >= 1656 AND x_counter <= 1661) OR (x_counter >= 1680 AND x_counter <= 1685) OR (x_counter >= 1689 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1703) OR (x_counter >= 1707 AND x_counter <= 1721)))
											OR	(y_counter = 423 AND ((x_counter >= 196 AND x_counter <= 201) OR (x_counter >= 205 AND x_counter <= 210) OR (x_counter >= 214 AND x_counter <= 219) OR (x_counter >= 223 AND x_counter <= 228) OR (x_counter >= 232 AND x_counter <= 237) OR (x_counter >= 241 AND x_counter <= 246) OR (x_counter >= 250 AND x_counter <= 255) OR (x_counter >= 259 AND x_counter <= 264) OR (x_counter >= 268 AND x_counter <= 273) OR (x_counter >= 286 AND x_counter <= 291) OR (x_counter >= 295 AND x_counter <= 300) OR (x_counter >= 304 AND x_counter <= 309) OR (x_counter >= 313 AND x_counter <= 318) OR (x_counter >= 322 AND x_counter <= 327) OR (x_counter >= 331 AND x_counter <= 336) OR (x_counter >= 340 AND x_counter <= 345) OR (x_counter >= 349 AND x_counter <= 354) OR (x_counter >= 358 AND x_counter <= 363) OR (x_counter >= 367 AND x_counter <= 372) OR (x_counter >= 376 AND x_counter <= 381) OR (x_counter >= 400 AND x_counter <= 405) OR (x_counter >= 409 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 423) OR (x_counter >= 427 AND x_counter <= 432) OR (x_counter >= 836 AND x_counter <= 841) OR (x_counter >= 845 AND x_counter <= 850) OR (x_counter >= 854 AND x_counter <= 859) OR (x_counter >= 863 AND x_counter <= 868) OR (x_counter >= 872 AND x_counter <= 877) OR (x_counter >= 881 AND x_counter <= 886) OR (x_counter >= 890 AND x_counter <= 895) OR (x_counter >= 899 AND x_counter <= 904) OR (x_counter >= 908 AND x_counter <= 913) OR (x_counter >= 926 AND x_counter <= 931) OR (x_counter >= 935 AND x_counter <= 940) OR (x_counter >= 944 AND x_counter <= 949) OR (x_counter >= 953 AND x_counter <= 958) OR (x_counter >= 962 AND x_counter <= 967) OR (x_counter >= 971 AND x_counter <= 976) OR (x_counter >= 980 AND x_counter <= 985) OR (x_counter >= 989 AND x_counter <= 994) OR (x_counter >= 998 AND x_counter <= 1003) OR (x_counter >= 1007 AND x_counter <= 1012) OR (x_counter >= 1016 AND x_counter <= 1021) OR (x_counter >= 1040 AND x_counter <= 1045) OR (x_counter >= 1049 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1063) OR (x_counter >= 1067 AND x_counter <= 1072) OR (x_counter >= 1476 AND x_counter <= 1481) OR (x_counter >= 1485 AND x_counter <= 1490) OR (x_counter >= 1494 AND x_counter <= 1499) OR (x_counter >= 1503 AND x_counter <= 1508) OR (x_counter >= 1512 AND x_counter <= 1517) OR (x_counter >= 1521 AND x_counter <= 1526) OR (x_counter >= 1530 AND x_counter <= 1535) OR (x_counter >= 1539 AND x_counter <= 1544) OR (x_counter >= 1548 AND x_counter <= 1553) OR (x_counter >= 1566 AND x_counter <= 1571) OR (x_counter >= 1575 AND x_counter <= 1580) OR (x_counter >= 1584 AND x_counter <= 1589) OR (x_counter >= 1593 AND x_counter <= 1598) OR (x_counter >= 1602 AND x_counter <= 1607) OR (x_counter >= 1611 AND x_counter <= 1616) OR (x_counter >= 1620 AND x_counter <= 1625) OR (x_counter >= 1629 AND x_counter <= 1634) OR (x_counter >= 1638 AND x_counter <= 1643) OR (x_counter >= 1647 AND x_counter <= 1652) OR (x_counter >= 1656 AND x_counter <= 1661) OR (x_counter >= 1680 AND x_counter <= 1685) OR (x_counter >= 1689 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1703) OR (x_counter >= 1707 AND x_counter <= 1712)))
											OR	(y_counter = 424 AND ((x_counter >= 196 AND x_counter <= 201) OR (x_counter >= 205 AND x_counter <= 210) OR (x_counter >= 214 AND x_counter <= 219) OR (x_counter >= 223 AND x_counter <= 228) OR (x_counter >= 232 AND x_counter <= 237) OR (x_counter >= 241 AND x_counter <= 246) OR (x_counter >= 250 AND x_counter <= 255) OR (x_counter >= 259 AND x_counter <= 264) OR (x_counter >= 268 AND x_counter <= 273) OR (x_counter >= 286 AND x_counter <= 291) OR (x_counter >= 295 AND x_counter <= 300) OR (x_counter >= 304 AND x_counter <= 309) OR (x_counter >= 313 AND x_counter <= 318) OR (x_counter >= 322 AND x_counter <= 327) OR (x_counter >= 331 AND x_counter <= 336) OR (x_counter >= 340 AND x_counter <= 345) OR (x_counter >= 349 AND x_counter <= 354) OR (x_counter >= 358 AND x_counter <= 363) OR (x_counter >= 367 AND x_counter <= 372) OR (x_counter >= 376 AND x_counter <= 381) OR (x_counter >= 400 AND x_counter <= 405) OR (x_counter >= 409 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 423) OR (x_counter >= 427 AND x_counter <= 432) OR (x_counter >= 836 AND x_counter <= 841) OR (x_counter >= 845 AND x_counter <= 850) OR (x_counter >= 854 AND x_counter <= 859) OR (x_counter >= 863 AND x_counter <= 868) OR (x_counter >= 872 AND x_counter <= 877) OR (x_counter >= 881 AND x_counter <= 886) OR (x_counter >= 890 AND x_counter <= 895) OR (x_counter >= 899 AND x_counter <= 904) OR (x_counter >= 908 AND x_counter <= 913) OR (x_counter >= 926 AND x_counter <= 931) OR (x_counter >= 935 AND x_counter <= 940) OR (x_counter >= 944 AND x_counter <= 949) OR (x_counter >= 953 AND x_counter <= 958) OR (x_counter >= 962 AND x_counter <= 967) OR (x_counter >= 971 AND x_counter <= 976) OR (x_counter >= 980 AND x_counter <= 985) OR (x_counter >= 989 AND x_counter <= 994) OR (x_counter >= 998 AND x_counter <= 1003) OR (x_counter >= 1007 AND x_counter <= 1012) OR (x_counter >= 1016 AND x_counter <= 1021) OR (x_counter >= 1040 AND x_counter <= 1045) OR (x_counter >= 1049 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1063) OR (x_counter >= 1067 AND x_counter <= 1072) OR (x_counter >= 1476 AND x_counter <= 1481) OR (x_counter >= 1485 AND x_counter <= 1490) OR (x_counter >= 1494 AND x_counter <= 1499) OR (x_counter >= 1503 AND x_counter <= 1508) OR (x_counter >= 1512 AND x_counter <= 1517) OR (x_counter >= 1521 AND x_counter <= 1526) OR (x_counter >= 1530 AND x_counter <= 1535) OR (x_counter >= 1539 AND x_counter <= 1544) OR (x_counter >= 1548 AND x_counter <= 1553) OR (x_counter >= 1566 AND x_counter <= 1571) OR (x_counter >= 1575 AND x_counter <= 1580) OR (x_counter >= 1584 AND x_counter <= 1589) OR (x_counter >= 1593 AND x_counter <= 1598) OR (x_counter >= 1602 AND x_counter <= 1607) OR (x_counter >= 1611 AND x_counter <= 1616) OR (x_counter >= 1620 AND x_counter <= 1625) OR (x_counter >= 1629 AND x_counter <= 1634) OR (x_counter >= 1638 AND x_counter <= 1643) OR (x_counter >= 1647 AND x_counter <= 1652) OR (x_counter >= 1656 AND x_counter <= 1661) OR (x_counter >= 1680 AND x_counter <= 1685) OR (x_counter >= 1689 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1703) OR (x_counter >= 1707 AND x_counter <= 1712)))
											OR	(y_counter = 425 AND ((x_counter >= 196 AND x_counter <= 201) OR (x_counter >= 205 AND x_counter <= 210) OR (x_counter >= 214 AND x_counter <= 219) OR (x_counter >= 223 AND x_counter <= 228) OR (x_counter >= 232 AND x_counter <= 237) OR (x_counter >= 241 AND x_counter <= 246) OR (x_counter >= 250 AND x_counter <= 255) OR (x_counter >= 259 AND x_counter <= 264) OR (x_counter >= 268 AND x_counter <= 273) OR (x_counter >= 286 AND x_counter <= 291) OR (x_counter >= 295 AND x_counter <= 300) OR (x_counter >= 304 AND x_counter <= 309) OR (x_counter >= 313 AND x_counter <= 318) OR (x_counter >= 322 AND x_counter <= 327) OR (x_counter >= 331 AND x_counter <= 336) OR (x_counter >= 340 AND x_counter <= 345) OR (x_counter >= 349 AND x_counter <= 354) OR (x_counter >= 358 AND x_counter <= 363) OR (x_counter >= 367 AND x_counter <= 372) OR (x_counter >= 376 AND x_counter <= 381) OR (x_counter >= 400 AND x_counter <= 405) OR (x_counter >= 409 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 423) OR (x_counter >= 427 AND x_counter <= 432) OR (x_counter >= 836 AND x_counter <= 841) OR (x_counter >= 845 AND x_counter <= 850) OR (x_counter >= 854 AND x_counter <= 859) OR (x_counter >= 863 AND x_counter <= 868) OR (x_counter >= 872 AND x_counter <= 877) OR (x_counter >= 881 AND x_counter <= 886) OR (x_counter >= 890 AND x_counter <= 895) OR (x_counter >= 899 AND x_counter <= 904) OR (x_counter >= 908 AND x_counter <= 913) OR (x_counter >= 926 AND x_counter <= 931) OR (x_counter >= 935 AND x_counter <= 940) OR (x_counter >= 944 AND x_counter <= 949) OR (x_counter >= 953 AND x_counter <= 958) OR (x_counter >= 962 AND x_counter <= 967) OR (x_counter >= 971 AND x_counter <= 976) OR (x_counter >= 980 AND x_counter <= 985) OR (x_counter >= 989 AND x_counter <= 994) OR (x_counter >= 998 AND x_counter <= 1003) OR (x_counter >= 1007 AND x_counter <= 1012) OR (x_counter >= 1016 AND x_counter <= 1021) OR (x_counter >= 1040 AND x_counter <= 1045) OR (x_counter >= 1049 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1063) OR (x_counter >= 1067 AND x_counter <= 1072) OR (x_counter >= 1476 AND x_counter <= 1481) OR (x_counter >= 1485 AND x_counter <= 1490) OR (x_counter >= 1494 AND x_counter <= 1499) OR (x_counter >= 1503 AND x_counter <= 1508) OR (x_counter >= 1512 AND x_counter <= 1517) OR (x_counter >= 1521 AND x_counter <= 1526) OR (x_counter >= 1530 AND x_counter <= 1535) OR (x_counter >= 1539 AND x_counter <= 1544) OR (x_counter >= 1548 AND x_counter <= 1553) OR (x_counter >= 1566 AND x_counter <= 1571) OR (x_counter >= 1575 AND x_counter <= 1580) OR (x_counter >= 1584 AND x_counter <= 1589) OR (x_counter >= 1593 AND x_counter <= 1598) OR (x_counter >= 1602 AND x_counter <= 1607) OR (x_counter >= 1611 AND x_counter <= 1616) OR (x_counter >= 1620 AND x_counter <= 1625) OR (x_counter >= 1629 AND x_counter <= 1634) OR (x_counter >= 1638 AND x_counter <= 1643) OR (x_counter >= 1647 AND x_counter <= 1652) OR (x_counter >= 1656 AND x_counter <= 1661) OR (x_counter >= 1680 AND x_counter <= 1685) OR (x_counter >= 1689 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1703) OR (x_counter >= 1707 AND x_counter <= 1712)))
											OR	(y_counter = 426 AND ((x_counter >= 196 AND x_counter <= 219) OR (x_counter >= 223 AND x_counter <= 246) OR (x_counter >= 250 AND x_counter <= 273) OR (x_counter >= 277 AND x_counter <= 282) OR (x_counter >= 286 AND x_counter <= 300) OR (x_counter >= 304 AND x_counter <= 309) OR (x_counter >= 313 AND x_counter <= 318) OR (x_counter >= 322 AND x_counter <= 336) OR (x_counter >= 340 AND x_counter <= 354) OR (x_counter >= 358 AND x_counter <= 372) OR (x_counter >= 376 AND x_counter <= 381) OR (x_counter >= 391 AND x_counter <= 396) OR (x_counter >= 400 AND x_counter <= 405) OR (x_counter >= 409 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 423) OR (x_counter >= 427 AND x_counter <= 441) OR (x_counter >= 836 AND x_counter <= 859) OR (x_counter >= 863 AND x_counter <= 886) OR (x_counter >= 890 AND x_counter <= 913) OR (x_counter >= 917 AND x_counter <= 922) OR (x_counter >= 926 AND x_counter <= 940) OR (x_counter >= 944 AND x_counter <= 949) OR (x_counter >= 953 AND x_counter <= 958) OR (x_counter >= 962 AND x_counter <= 976) OR (x_counter >= 980 AND x_counter <= 994) OR (x_counter >= 998 AND x_counter <= 1012) OR (x_counter >= 1016 AND x_counter <= 1021) OR (x_counter >= 1031 AND x_counter <= 1036) OR (x_counter >= 1040 AND x_counter <= 1045) OR (x_counter >= 1049 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1063) OR (x_counter >= 1067 AND x_counter <= 1081) OR (x_counter >= 1476 AND x_counter <= 1499) OR (x_counter >= 1503 AND x_counter <= 1526) OR (x_counter >= 1530 AND x_counter <= 1553) OR (x_counter >= 1557 AND x_counter <= 1562) OR (x_counter >= 1566 AND x_counter <= 1580) OR (x_counter >= 1584 AND x_counter <= 1589) OR (x_counter >= 1593 AND x_counter <= 1598) OR (x_counter >= 1602 AND x_counter <= 1616) OR (x_counter >= 1620 AND x_counter <= 1634) OR (x_counter >= 1638 AND x_counter <= 1652) OR (x_counter >= 1656 AND x_counter <= 1661) OR (x_counter >= 1671 AND x_counter <= 1676) OR (x_counter >= 1680 AND x_counter <= 1685) OR (x_counter >= 1689 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1703) OR (x_counter >= 1707 AND x_counter <= 1721)))
											OR	(y_counter = 427 AND ((x_counter >= 196 AND x_counter <= 219) OR (x_counter >= 223 AND x_counter <= 246) OR (x_counter >= 250 AND x_counter <= 273) OR (x_counter >= 277 AND x_counter <= 282) OR (x_counter >= 286 AND x_counter <= 300) OR (x_counter >= 304 AND x_counter <= 309) OR (x_counter >= 313 AND x_counter <= 318) OR (x_counter >= 322 AND x_counter <= 336) OR (x_counter >= 340 AND x_counter <= 354) OR (x_counter >= 358 AND x_counter <= 372) OR (x_counter >= 376 AND x_counter <= 381) OR (x_counter >= 391 AND x_counter <= 396) OR (x_counter >= 400 AND x_counter <= 405) OR (x_counter >= 409 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 423) OR (x_counter >= 427 AND x_counter <= 441) OR (x_counter >= 836 AND x_counter <= 859) OR (x_counter >= 863 AND x_counter <= 886) OR (x_counter >= 890 AND x_counter <= 913) OR (x_counter >= 917 AND x_counter <= 922) OR (x_counter >= 926 AND x_counter <= 940) OR (x_counter >= 944 AND x_counter <= 949) OR (x_counter >= 953 AND x_counter <= 958) OR (x_counter >= 962 AND x_counter <= 976) OR (x_counter >= 980 AND x_counter <= 994) OR (x_counter >= 998 AND x_counter <= 1012) OR (x_counter >= 1016 AND x_counter <= 1021) OR (x_counter >= 1031 AND x_counter <= 1036) OR (x_counter >= 1040 AND x_counter <= 1045) OR (x_counter >= 1049 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1063) OR (x_counter >= 1067 AND x_counter <= 1081) OR (x_counter >= 1476 AND x_counter <= 1499) OR (x_counter >= 1503 AND x_counter <= 1526) OR (x_counter >= 1530 AND x_counter <= 1553) OR (x_counter >= 1557 AND x_counter <= 1562) OR (x_counter >= 1566 AND x_counter <= 1580) OR (x_counter >= 1584 AND x_counter <= 1589) OR (x_counter >= 1593 AND x_counter <= 1598) OR (x_counter >= 1602 AND x_counter <= 1616) OR (x_counter >= 1620 AND x_counter <= 1634) OR (x_counter >= 1638 AND x_counter <= 1652) OR (x_counter >= 1656 AND x_counter <= 1661) OR (x_counter >= 1671 AND x_counter <= 1676) OR (x_counter >= 1680 AND x_counter <= 1685) OR (x_counter >= 1689 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1703) OR (x_counter >= 1707 AND x_counter <= 1721)))
											OR	(y_counter = 428 AND ((x_counter >= 196 AND x_counter <= 219) OR (x_counter >= 223 AND x_counter <= 246) OR (x_counter >= 250 AND x_counter <= 273) OR (x_counter >= 277 AND x_counter <= 282) OR (x_counter >= 286 AND x_counter <= 300) OR (x_counter >= 304 AND x_counter <= 309) OR (x_counter >= 313 AND x_counter <= 318) OR (x_counter >= 322 AND x_counter <= 336) OR (x_counter >= 340 AND x_counter <= 354) OR (x_counter >= 358 AND x_counter <= 372) OR (x_counter >= 376 AND x_counter <= 381) OR (x_counter >= 391 AND x_counter <= 396) OR (x_counter >= 400 AND x_counter <= 405) OR (x_counter >= 409 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 423) OR (x_counter >= 427 AND x_counter <= 441) OR (x_counter >= 836 AND x_counter <= 859) OR (x_counter >= 863 AND x_counter <= 886) OR (x_counter >= 890 AND x_counter <= 913) OR (x_counter >= 917 AND x_counter <= 922) OR (x_counter >= 926 AND x_counter <= 940) OR (x_counter >= 944 AND x_counter <= 949) OR (x_counter >= 953 AND x_counter <= 958) OR (x_counter >= 962 AND x_counter <= 976) OR (x_counter >= 980 AND x_counter <= 994) OR (x_counter >= 998 AND x_counter <= 1012) OR (x_counter >= 1016 AND x_counter <= 1021) OR (x_counter >= 1031 AND x_counter <= 1036) OR (x_counter >= 1040 AND x_counter <= 1045) OR (x_counter >= 1049 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1063) OR (x_counter >= 1067 AND x_counter <= 1081) OR (x_counter >= 1476 AND x_counter <= 1499) OR (x_counter >= 1503 AND x_counter <= 1526) OR (x_counter >= 1530 AND x_counter <= 1553) OR (x_counter >= 1557 AND x_counter <= 1562) OR (x_counter >= 1566 AND x_counter <= 1580) OR (x_counter >= 1584 AND x_counter <= 1589) OR (x_counter >= 1593 AND x_counter <= 1598) OR (x_counter >= 1602 AND x_counter <= 1616) OR (x_counter >= 1620 AND x_counter <= 1634) OR (x_counter >= 1638 AND x_counter <= 1652) OR (x_counter >= 1656 AND x_counter <= 1661) OR (x_counter >= 1671 AND x_counter <= 1676) OR (x_counter >= 1680 AND x_counter <= 1685) OR (x_counter >= 1689 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1703) OR (x_counter >= 1707 AND x_counter <= 1721)))
											OR	(y_counter = 429 AND ((x_counter >= 196 AND x_counter <= 219) OR (x_counter >= 223 AND x_counter <= 246) OR (x_counter >= 250 AND x_counter <= 273) OR (x_counter >= 277 AND x_counter <= 282) OR (x_counter >= 286 AND x_counter <= 300) OR (x_counter >= 304 AND x_counter <= 309) OR (x_counter >= 313 AND x_counter <= 318) OR (x_counter >= 322 AND x_counter <= 336) OR (x_counter >= 340 AND x_counter <= 354) OR (x_counter >= 358 AND x_counter <= 372) OR (x_counter >= 376 AND x_counter <= 381) OR (x_counter >= 391 AND x_counter <= 396) OR (x_counter >= 400 AND x_counter <= 405) OR (x_counter >= 409 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 423) OR (x_counter >= 427 AND x_counter <= 441) OR (x_counter >= 836 AND x_counter <= 859) OR (x_counter >= 863 AND x_counter <= 886) OR (x_counter >= 890 AND x_counter <= 913) OR (x_counter >= 917 AND x_counter <= 922) OR (x_counter >= 926 AND x_counter <= 940) OR (x_counter >= 944 AND x_counter <= 949) OR (x_counter >= 953 AND x_counter <= 958) OR (x_counter >= 962 AND x_counter <= 976) OR (x_counter >= 980 AND x_counter <= 994) OR (x_counter >= 998 AND x_counter <= 1012) OR (x_counter >= 1016 AND x_counter <= 1021) OR (x_counter >= 1031 AND x_counter <= 1036) OR (x_counter >= 1040 AND x_counter <= 1045) OR (x_counter >= 1049 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1063) OR (x_counter >= 1067 AND x_counter <= 1081) OR (x_counter >= 1476 AND x_counter <= 1499) OR (x_counter >= 1503 AND x_counter <= 1526) OR (x_counter >= 1530 AND x_counter <= 1553) OR (x_counter >= 1557 AND x_counter <= 1562) OR (x_counter >= 1566 AND x_counter <= 1580) OR (x_counter >= 1584 AND x_counter <= 1589) OR (x_counter >= 1593 AND x_counter <= 1598) OR (x_counter >= 1602 AND x_counter <= 1616) OR (x_counter >= 1620 AND x_counter <= 1634) OR (x_counter >= 1638 AND x_counter <= 1652) OR (x_counter >= 1656 AND x_counter <= 1661) OR (x_counter >= 1671 AND x_counter <= 1676) OR (x_counter >= 1680 AND x_counter <= 1685) OR (x_counter >= 1689 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1703) OR (x_counter >= 1707 AND x_counter <= 1721)))
											OR	(y_counter = 430 AND ((x_counter >= 196 AND x_counter <= 219) OR (x_counter >= 223 AND x_counter <= 246) OR (x_counter >= 250 AND x_counter <= 273) OR (x_counter >= 277 AND x_counter <= 282) OR (x_counter >= 286 AND x_counter <= 300) OR (x_counter >= 304 AND x_counter <= 309) OR (x_counter >= 313 AND x_counter <= 318) OR (x_counter >= 322 AND x_counter <= 336) OR (x_counter >= 340 AND x_counter <= 354) OR (x_counter >= 358 AND x_counter <= 372) OR (x_counter >= 376 AND x_counter <= 381) OR (x_counter >= 391 AND x_counter <= 396) OR (x_counter >= 400 AND x_counter <= 405) OR (x_counter >= 409 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 423) OR (x_counter >= 427 AND x_counter <= 441) OR (x_counter >= 836 AND x_counter <= 859) OR (x_counter >= 863 AND x_counter <= 886) OR (x_counter >= 890 AND x_counter <= 913) OR (x_counter >= 917 AND x_counter <= 922) OR (x_counter >= 926 AND x_counter <= 940) OR (x_counter >= 944 AND x_counter <= 949) OR (x_counter >= 953 AND x_counter <= 958) OR (x_counter >= 962 AND x_counter <= 976) OR (x_counter >= 980 AND x_counter <= 994) OR (x_counter >= 998 AND x_counter <= 1012) OR (x_counter >= 1016 AND x_counter <= 1021) OR (x_counter >= 1031 AND x_counter <= 1036) OR (x_counter >= 1040 AND x_counter <= 1045) OR (x_counter >= 1049 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1063) OR (x_counter >= 1067 AND x_counter <= 1081) OR (x_counter >= 1476 AND x_counter <= 1499) OR (x_counter >= 1503 AND x_counter <= 1526) OR (x_counter >= 1530 AND x_counter <= 1553) OR (x_counter >= 1557 AND x_counter <= 1562) OR (x_counter >= 1566 AND x_counter <= 1580) OR (x_counter >= 1584 AND x_counter <= 1589) OR (x_counter >= 1593 AND x_counter <= 1598) OR (x_counter >= 1602 AND x_counter <= 1616) OR (x_counter >= 1620 AND x_counter <= 1634) OR (x_counter >= 1638 AND x_counter <= 1652) OR (x_counter >= 1656 AND x_counter <= 1661) OR (x_counter >= 1671 AND x_counter <= 1676) OR (x_counter >= 1680 AND x_counter <= 1685) OR (x_counter >= 1689 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1703) OR (x_counter >= 1707 AND x_counter <= 1721)))
											OR	(y_counter = 431 AND ((x_counter >= 196 AND x_counter <= 219) OR (x_counter >= 223 AND x_counter <= 246) OR (x_counter >= 250 AND x_counter <= 273) OR (x_counter >= 277 AND x_counter <= 282) OR (x_counter >= 286 AND x_counter <= 300) OR (x_counter >= 304 AND x_counter <= 309) OR (x_counter >= 313 AND x_counter <= 318) OR (x_counter >= 322 AND x_counter <= 336) OR (x_counter >= 340 AND x_counter <= 354) OR (x_counter >= 358 AND x_counter <= 372) OR (x_counter >= 376 AND x_counter <= 381) OR (x_counter >= 391 AND x_counter <= 396) OR (x_counter >= 400 AND x_counter <= 405) OR (x_counter >= 409 AND x_counter <= 414) OR (x_counter >= 418 AND x_counter <= 423) OR (x_counter >= 427 AND x_counter <= 441) OR (x_counter >= 836 AND x_counter <= 859) OR (x_counter >= 863 AND x_counter <= 886) OR (x_counter >= 890 AND x_counter <= 913) OR (x_counter >= 917 AND x_counter <= 922) OR (x_counter >= 926 AND x_counter <= 940) OR (x_counter >= 944 AND x_counter <= 949) OR (x_counter >= 953 AND x_counter <= 958) OR (x_counter >= 962 AND x_counter <= 976) OR (x_counter >= 980 AND x_counter <= 994) OR (x_counter >= 998 AND x_counter <= 1012) OR (x_counter >= 1016 AND x_counter <= 1021) OR (x_counter >= 1031 AND x_counter <= 1036) OR (x_counter >= 1040 AND x_counter <= 1045) OR (x_counter >= 1049 AND x_counter <= 1054) OR (x_counter >= 1058 AND x_counter <= 1063) OR (x_counter >= 1067 AND x_counter <= 1081) OR (x_counter >= 1476 AND x_counter <= 1499) OR (x_counter >= 1503 AND x_counter <= 1526) OR (x_counter >= 1530 AND x_counter <= 1553) OR (x_counter >= 1557 AND x_counter <= 1562) OR (x_counter >= 1566 AND x_counter <= 1580) OR (x_counter >= 1584 AND x_counter <= 1589) OR (x_counter >= 1593 AND x_counter <= 1598) OR (x_counter >= 1602 AND x_counter <= 1616) OR (x_counter >= 1620 AND x_counter <= 1634) OR (x_counter >= 1638 AND x_counter <= 1652) OR (x_counter >= 1656 AND x_counter <= 1661) OR (x_counter >= 1671 AND x_counter <= 1676) OR (x_counter >= 1680 AND x_counter <= 1685) OR (x_counter >= 1689 AND x_counter <= 1694) OR (x_counter >= 1698 AND x_counter <= 1703) OR (x_counter >= 1707 AND x_counter <= 1721)))
											OR	(y_counter = 432 AND ((x_counter >= 322 AND x_counter <= 327) OR (x_counter >= 962 AND x_counter <= 967) OR (x_counter >= 1602 AND x_counter <= 1607)))
											OR	(y_counter = 433 AND ((x_counter >= 322 AND x_counter <= 327) OR (x_counter >= 962 AND x_counter <= 967) OR (x_counter >= 1602 AND x_counter <= 1607)))
											OR	(y_counter = 434 AND ((x_counter >= 322 AND x_counter <= 327) OR (x_counter >= 962 AND x_counter <= 967) OR (x_counter >= 1602 AND x_counter <= 1607)))
											OR	(y_counter = 435 AND ((x_counter >= 322 AND x_counter <= 327) OR (x_counter >= 962 AND x_counter <= 967) OR (x_counter >= 1602 AND x_counter <= 1607)))
											OR	(y_counter = 436 AND ((x_counter >= 322 AND x_counter <= 327) OR (x_counter >= 962 AND x_counter <= 967) OR (x_counter >= 1602 AND x_counter <= 1607)))
											OR	(y_counter = 437 AND ((x_counter >= 322 AND x_counter <= 327) OR (x_counter >= 962 AND x_counter <= 967) OR (x_counter >= 1602 AND x_counter <= 1607)))
											OR	(y_counter = 438 AND ((x_counter >= 322 AND x_counter <= 327) OR (x_counter >= 962 AND x_counter <= 967) OR (x_counter >= 1602 AND x_counter <= 1607)))
											OR	(y_counter = 439 AND ((x_counter >= 322 AND x_counter <= 327) OR (x_counter >= 962 AND x_counter <= 967) OR (x_counter >= 1602 AND x_counter <= 1607)))
											OR	(y_counter = 440 AND ((x_counter >= 322 AND x_counter <= 327) OR (x_counter >= 962 AND x_counter <= 967) OR (x_counter >= 1602 AND x_counter <= 1607)))
											else "000";


end Behavioral;

