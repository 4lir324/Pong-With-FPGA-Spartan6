
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity gameover_menu is
--FPGA pin decleration
    Port (		 clk			 :		in std_logic;
					 reset 		 :		in std_logic;
					 x_counter   :  	in integer range 0 to 640;
                y_counter   :   	in integer range 0 to 480;
                RGB         :   	out STD_LOGIC_VECTOR(2 downto 0));  --VGA RGB output
end gameover_menu;

architecture Behavioral of gameover_menu is

    signal animation_on : std_logic; --flashing the "PRESS ANY KEY"
begin

-------------------------------------------Animation-----------------------------------------------------
    process(clk,reset)
        variable    animation_timer_var : integer range 0 to 25000000;
        begin
            if(reset = '1') then
                animation_timer_var := 0;
                animation_on <= '0';
                
            elsif (clk'event and clk = '1') then
                animation_timer_var := animation_timer_var + 1;
                    if(animation_timer_var = 25000000) then
                        animation_timer_var := 0;
                        animation_on <= not(animation_on);
                    end if;
            end if;
        
        end process;

				RGB   <= "111" when		       ( y_counter = 169 AND ((x_counter >= 181 AND x_counter <= 198 ) OR (x_counter >= 346 AND x_counter <= 363 )))
                                        OR ( y_counter = 170 AND ((x_counter >= 181 AND x_counter <= 198 ) OR (x_counter >= 346 AND x_counter <= 363 )))
                                        OR ( y_counter = 171 AND ((x_counter >= 181 AND x_counter <= 198 ) OR (x_counter >= 346 AND x_counter <= 363 )))
                                        OR ( y_counter = 172 AND ((x_counter >= 181 AND x_counter <= 198 ) OR (x_counter >= 346 AND x_counter <= 363 )))
                                        OR ( y_counter = 173 AND ((x_counter >= 177 AND x_counter <= 186 ) OR (x_counter >= 193 AND x_counter <= 202 ) OR (x_counter >= 342 AND x_counter <= 351 ) OR (x_counter >= 358 AND x_counter <= 367 )))
                                        OR ( y_counter = 174 AND ((x_counter >= 177 AND x_counter <= 186 ) OR (x_counter >= 193 AND x_counter <= 202 ) OR (x_counter >= 342 AND x_counter <= 351 ) OR (x_counter >= 358 AND x_counter <= 367 )))
                                        OR ( y_counter = 175 AND ((x_counter >= 177 AND x_counter <= 186 ) OR (x_counter >= 193 AND x_counter <= 202 ) OR (x_counter >= 342 AND x_counter <= 351 ) OR (x_counter >= 358 AND x_counter <= 367 )))
                                        OR ( y_counter = 176 AND ((x_counter >= 177 AND x_counter <= 186 ) OR (x_counter >= 193 AND x_counter <= 202 ) OR (x_counter >= 342 AND x_counter <= 351 ) OR (x_counter >= 358 AND x_counter <= 367 )))
                                        OR ( y_counter = 177 AND ((x_counter >= 177 AND x_counter <= 186 ) OR (x_counter >= 193 AND x_counter <= 202 ) OR (x_counter >= 214 AND x_counter <= 231 ) OR (x_counter >= 243 AND x_counter <= 268 ) OR (x_counter >= 280 AND x_counter <= 297 ) OR (x_counter >= 342 AND x_counter <= 351 ) OR (x_counter >= 358 AND x_counter <= 367 ) OR (x_counter >= 375 AND x_counter <= 384 ) OR (x_counter >= 391 AND x_counter <= 400 ) OR (x_counter >= 412 AND x_counter <= 429 ) OR (x_counter >= 441 AND x_counter <= 450 ) OR (x_counter >= 457 AND x_counter <= 466 )))
                                        OR ( y_counter = 178 AND ((x_counter >= 177 AND x_counter <= 186 ) OR (x_counter >= 193 AND x_counter <= 202 ) OR (x_counter >= 214 AND x_counter <= 231 ) OR (x_counter >= 243 AND x_counter <= 268 ) OR (x_counter >= 280 AND x_counter <= 297 ) OR (x_counter >= 342 AND x_counter <= 351 ) OR (x_counter >= 358 AND x_counter <= 367 ) OR (x_counter >= 375 AND x_counter <= 384 ) OR (x_counter >= 391 AND x_counter <= 400 ) OR (x_counter >= 412 AND x_counter <= 429 ) OR (x_counter >= 441 AND x_counter <= 450 ) OR (x_counter >= 457 AND x_counter <= 466 )))
                                        OR ( y_counter = 179 AND ((x_counter >= 177 AND x_counter <= 186 ) OR (x_counter >= 193 AND x_counter <= 202 ) OR (x_counter >= 214 AND x_counter <= 231 ) OR (x_counter >= 243 AND x_counter <= 268 ) OR (x_counter >= 280 AND x_counter <= 297 ) OR (x_counter >= 342 AND x_counter <= 351 ) OR (x_counter >= 358 AND x_counter <= 367 ) OR (x_counter >= 375 AND x_counter <= 384 ) OR (x_counter >= 391 AND x_counter <= 400 ) OR (x_counter >= 412 AND x_counter <= 429 ) OR (x_counter >= 441 AND x_counter <= 450 ) OR (x_counter >= 457 AND x_counter <= 466 )))
                                        OR ( y_counter = 180 AND ((x_counter >= 177 AND x_counter <= 186 ) OR (x_counter >= 193 AND x_counter <= 202 ) OR (x_counter >= 214 AND x_counter <= 231 ) OR (x_counter >= 243 AND x_counter <= 268 ) OR (x_counter >= 280 AND x_counter <= 297 ) OR (x_counter >= 342 AND x_counter <= 351 ) OR (x_counter >= 358 AND x_counter <= 367 ) OR (x_counter >= 375 AND x_counter <= 384 ) OR (x_counter >= 391 AND x_counter <= 400 ) OR (x_counter >= 412 AND x_counter <= 429 ) OR (x_counter >= 441 AND x_counter <= 450 ) OR (x_counter >= 457 AND x_counter <= 466 )))
                                        OR ( y_counter = 181 AND ((x_counter >= 177 AND x_counter <= 186 ) OR (x_counter >= 226 AND x_counter <= 235 ) OR (x_counter >= 243 AND x_counter <= 252 ) OR (x_counter >= 255 AND x_counter <= 260 ) OR (x_counter >= 263 AND x_counter <= 272 ) OR (x_counter >= 276 AND x_counter <= 285 ) OR (x_counter >= 292 AND x_counter <= 301 ) OR (x_counter >= 342 AND x_counter <= 351 ) OR (x_counter >= 358 AND x_counter <= 367 ) OR (x_counter >= 375 AND x_counter <= 384 ) OR (x_counter >= 391 AND x_counter <= 400 ) OR (x_counter >= 408 AND x_counter <= 417 ) OR (x_counter >= 424 AND x_counter <= 433 ) OR (x_counter >= 441 AND x_counter <= 450 ) OR (x_counter >= 453 AND x_counter <= 466 )))
                                        OR ( y_counter = 182 AND ((x_counter >= 177 AND x_counter <= 186 ) OR (x_counter >= 226 AND x_counter <= 235 ) OR (x_counter >= 243 AND x_counter <= 252 ) OR (x_counter >= 255 AND x_counter <= 260 ) OR (x_counter >= 263 AND x_counter <= 272 ) OR (x_counter >= 276 AND x_counter <= 285 ) OR (x_counter >= 292 AND x_counter <= 301 ) OR (x_counter >= 342 AND x_counter <= 351 ) OR (x_counter >= 358 AND x_counter <= 367 ) OR (x_counter >= 375 AND x_counter <= 384 ) OR (x_counter >= 391 AND x_counter <= 400 ) OR (x_counter >= 408 AND x_counter <= 417 ) OR (x_counter >= 424 AND x_counter <= 433 ) OR (x_counter >= 441 AND x_counter <= 450 ) OR (x_counter >= 453 AND x_counter <= 466 )))
                                        OR ( y_counter = 183 AND ((x_counter >= 177 AND x_counter <= 186 ) OR (x_counter >= 226 AND x_counter <= 235 ) OR (x_counter >= 243 AND x_counter <= 252 ) OR (x_counter >= 255 AND x_counter <= 260 ) OR (x_counter >= 263 AND x_counter <= 272 ) OR (x_counter >= 276 AND x_counter <= 285 ) OR (x_counter >= 292 AND x_counter <= 301 ) OR (x_counter >= 342 AND x_counter <= 351 ) OR (x_counter >= 358 AND x_counter <= 367 ) OR (x_counter >= 375 AND x_counter <= 384 ) OR (x_counter >= 391 AND x_counter <= 400 ) OR (x_counter >= 408 AND x_counter <= 417 ) OR (x_counter >= 424 AND x_counter <= 433 ) OR (x_counter >= 441 AND x_counter <= 450 ) OR (x_counter >= 453 AND x_counter <= 466 )))
                                        OR ( y_counter = 184 AND ((x_counter >= 177 AND x_counter <= 186 ) OR (x_counter >= 226 AND x_counter <= 235 ) OR (x_counter >= 243 AND x_counter <= 252 ) OR (x_counter >= 255 AND x_counter <= 260 ) OR (x_counter >= 263 AND x_counter <= 272 ) OR (x_counter >= 276 AND x_counter <= 285 ) OR (x_counter >= 292 AND x_counter <= 301 ) OR (x_counter >= 342 AND x_counter <= 351 ) OR (x_counter >= 358 AND x_counter <= 367 ) OR (x_counter >= 375 AND x_counter <= 384 ) OR (x_counter >= 391 AND x_counter <= 400 ) OR (x_counter >= 408 AND x_counter <= 417 ) OR (x_counter >= 424 AND x_counter <= 433 ) OR (x_counter >= 441 AND x_counter <= 450 ) OR (x_counter >= 453 AND x_counter <= 466 )))
                                        OR ( y_counter = 185 AND ((x_counter >= 177 AND x_counter <= 186 ) OR (x_counter >= 226 AND x_counter <= 235 ) OR (x_counter >= 243 AND x_counter <= 252 ) OR (x_counter >= 255 AND x_counter <= 260 ) OR (x_counter >= 263 AND x_counter <= 272 ) OR (x_counter >= 276 AND x_counter <= 285 ) OR (x_counter >= 292 AND x_counter <= 301 ) OR (x_counter >= 342 AND x_counter <= 351 ) OR (x_counter >= 358 AND x_counter <= 367 ) OR (x_counter >= 375 AND x_counter <= 384 ) OR (x_counter >= 391 AND x_counter <= 400 ) OR (x_counter >= 408 AND x_counter <= 417 ) OR (x_counter >= 424 AND x_counter <= 433 ) OR (x_counter >= 441 AND x_counter <= 454 )))
                                        OR ( y_counter = 186 AND ((x_counter >= 177 AND x_counter <= 186 ) OR (x_counter >= 226 AND x_counter <= 235 ) OR (x_counter >= 243 AND x_counter <= 252 ) OR (x_counter >= 255 AND x_counter <= 260 ) OR (x_counter >= 263 AND x_counter <= 272 ) OR (x_counter >= 276 AND x_counter <= 285 ) OR (x_counter >= 292 AND x_counter <= 301 ) OR (x_counter >= 342 AND x_counter <= 351 ) OR (x_counter >= 358 AND x_counter <= 367 ) OR (x_counter >= 375 AND x_counter <= 384 ) OR (x_counter >= 391 AND x_counter <= 400 ) OR (x_counter >= 408 AND x_counter <= 417 ) OR (x_counter >= 424 AND x_counter <= 433 ) OR (x_counter >= 441 AND x_counter <= 454 )))
                                        OR ( y_counter = 187 AND ((x_counter >= 177 AND x_counter <= 186 ) OR (x_counter >= 226 AND x_counter <= 235 ) OR (x_counter >= 243 AND x_counter <= 252 ) OR (x_counter >= 255 AND x_counter <= 260 ) OR (x_counter >= 263 AND x_counter <= 272 ) OR (x_counter >= 276 AND x_counter <= 285 ) OR (x_counter >= 292 AND x_counter <= 301 ) OR (x_counter >= 342 AND x_counter <= 351 ) OR (x_counter >= 358 AND x_counter <= 367 ) OR (x_counter >= 375 AND x_counter <= 384 ) OR (x_counter >= 391 AND x_counter <= 400 ) OR (x_counter >= 408 AND x_counter <= 417 ) OR (x_counter >= 424 AND x_counter <= 433 ) OR (x_counter >= 441 AND x_counter <= 454 )))
                                        OR ( y_counter = 188 AND ((x_counter >= 177 AND x_counter <= 186 ) OR (x_counter >= 226 AND x_counter <= 235 ) OR (x_counter >= 243 AND x_counter <= 252 ) OR (x_counter >= 255 AND x_counter <= 260 ) OR (x_counter >= 263 AND x_counter <= 272 ) OR (x_counter >= 276 AND x_counter <= 285 ) OR (x_counter >= 292 AND x_counter <= 301 ) OR (x_counter >= 342 AND x_counter <= 351 ) OR (x_counter >= 358 AND x_counter <= 367 ) OR (x_counter >= 375 AND x_counter <= 384 ) OR (x_counter >= 391 AND x_counter <= 400 ) OR (x_counter >= 408 AND x_counter <= 417 ) OR (x_counter >= 424 AND x_counter <= 433 ) OR (x_counter >= 441 AND x_counter <= 454 )))
                                        OR ( y_counter = 189 AND ((x_counter >= 177 AND x_counter <= 186 ) OR (x_counter >= 189 AND x_counter <= 202 ) OR (x_counter >= 214 AND x_counter <= 235 ) OR (x_counter >= 243 AND x_counter <= 252 ) OR (x_counter >= 255 AND x_counter <= 260 ) OR (x_counter >= 263 AND x_counter <= 272 ) OR (x_counter >= 276 AND x_counter <= 301 ) OR (x_counter >= 342 AND x_counter <= 351 ) OR (x_counter >= 358 AND x_counter <= 367 ) OR (x_counter >= 375 AND x_counter <= 384 ) OR (x_counter >= 391 AND x_counter <= 400 ) OR (x_counter >= 408 AND x_counter <= 433 ) OR (x_counter >= 441 AND x_counter <= 450 )))
                                        OR ( y_counter = 190 AND ((x_counter >= 177 AND x_counter <= 186 ) OR (x_counter >= 189 AND x_counter <= 202 ) OR (x_counter >= 214 AND x_counter <= 235 ) OR (x_counter >= 243 AND x_counter <= 252 ) OR (x_counter >= 255 AND x_counter <= 260 ) OR (x_counter >= 263 AND x_counter <= 272 ) OR (x_counter >= 276 AND x_counter <= 301 ) OR (x_counter >= 342 AND x_counter <= 351 ) OR (x_counter >= 358 AND x_counter <= 367 ) OR (x_counter >= 375 AND x_counter <= 384 ) OR (x_counter >= 391 AND x_counter <= 400 ) OR (x_counter >= 408 AND x_counter <= 433 ) OR (x_counter >= 441 AND x_counter <= 450 )))
                                        OR ( y_counter = 191 AND ((x_counter >= 177 AND x_counter <= 186 ) OR (x_counter >= 189 AND x_counter <= 202 ) OR (x_counter >= 214 AND x_counter <= 235 ) OR (x_counter >= 243 AND x_counter <= 252 ) OR (x_counter >= 255 AND x_counter <= 260 ) OR (x_counter >= 263 AND x_counter <= 272 ) OR (x_counter >= 276 AND x_counter <= 301 ) OR (x_counter >= 342 AND x_counter <= 351 ) OR (x_counter >= 358 AND x_counter <= 367 ) OR (x_counter >= 375 AND x_counter <= 384 ) OR (x_counter >= 391 AND x_counter <= 400 ) OR (x_counter >= 408 AND x_counter <= 433 ) OR (x_counter >= 441 AND x_counter <= 450 )))
                                        OR ( y_counter = 192 AND ((x_counter >= 177 AND x_counter <= 186 ) OR (x_counter >= 189 AND x_counter <= 202 ) OR (x_counter >= 214 AND x_counter <= 235 ) OR (x_counter >= 243 AND x_counter <= 252 ) OR (x_counter >= 255 AND x_counter <= 260 ) OR (x_counter >= 263 AND x_counter <= 272 ) OR (x_counter >= 276 AND x_counter <= 301 ) OR (x_counter >= 342 AND x_counter <= 351 ) OR (x_counter >= 358 AND x_counter <= 367 ) OR (x_counter >= 375 AND x_counter <= 384 ) OR (x_counter >= 391 AND x_counter <= 400 ) OR (x_counter >= 408 AND x_counter <= 433 ) OR (x_counter >= 441 AND x_counter <= 450 )))
                                        OR ( y_counter = 193 AND ((x_counter >= 177 AND x_counter <= 186 ) OR (x_counter >= 193 AND x_counter <= 202 ) OR (x_counter >= 210 AND x_counter <= 219 ) OR (x_counter >= 226 AND x_counter <= 235 ) OR (x_counter >= 243 AND x_counter <= 252 ) OR (x_counter >= 255 AND x_counter <= 260 ) OR (x_counter >= 263 AND x_counter <= 272 ) OR (x_counter >= 276 AND x_counter <= 285 ) OR (x_counter >= 342 AND x_counter <= 351 ) OR (x_counter >= 358 AND x_counter <= 367 ) OR (x_counter >= 375 AND x_counter <= 384 ) OR (x_counter >= 391 AND x_counter <= 400 ) OR (x_counter >= 408 AND x_counter <= 417 ) OR (x_counter >= 441 AND x_counter <= 450 )))
                                        OR ( y_counter = 194 AND ((x_counter >= 177 AND x_counter <= 186 ) OR (x_counter >= 193 AND x_counter <= 202 ) OR (x_counter >= 210 AND x_counter <= 219 ) OR (x_counter >= 226 AND x_counter <= 235 ) OR (x_counter >= 243 AND x_counter <= 252 ) OR (x_counter >= 255 AND x_counter <= 260 ) OR (x_counter >= 263 AND x_counter <= 272 ) OR (x_counter >= 276 AND x_counter <= 285 ) OR (x_counter >= 342 AND x_counter <= 351 ) OR (x_counter >= 358 AND x_counter <= 367 ) OR (x_counter >= 375 AND x_counter <= 384 ) OR (x_counter >= 391 AND x_counter <= 400 ) OR (x_counter >= 408 AND x_counter <= 417 ) OR (x_counter >= 441 AND x_counter <= 450 )))
                                        OR ( y_counter = 195 AND ((x_counter >= 177 AND x_counter <= 186 ) OR (x_counter >= 193 AND x_counter <= 202 ) OR (x_counter >= 210 AND x_counter <= 219 ) OR (x_counter >= 226 AND x_counter <= 235 ) OR (x_counter >= 243 AND x_counter <= 252 ) OR (x_counter >= 255 AND x_counter <= 260 ) OR (x_counter >= 263 AND x_counter <= 272 ) OR (x_counter >= 276 AND x_counter <= 285 ) OR (x_counter >= 342 AND x_counter <= 351 ) OR (x_counter >= 358 AND x_counter <= 367 ) OR (x_counter >= 375 AND x_counter <= 384 ) OR (x_counter >= 391 AND x_counter <= 400 ) OR (x_counter >= 408 AND x_counter <= 417 ) OR (x_counter >= 441 AND x_counter <= 450 )))
                                        OR ( y_counter = 196 AND ((x_counter >= 177 AND x_counter <= 186 ) OR (x_counter >= 193 AND x_counter <= 202 ) OR (x_counter >= 210 AND x_counter <= 219 ) OR (x_counter >= 226 AND x_counter <= 235 ) OR (x_counter >= 243 AND x_counter <= 252 ) OR (x_counter >= 255 AND x_counter <= 260 ) OR (x_counter >= 263 AND x_counter <= 272 ) OR (x_counter >= 276 AND x_counter <= 285 ) OR (x_counter >= 342 AND x_counter <= 351 ) OR (x_counter >= 358 AND x_counter <= 367 ) OR (x_counter >= 375 AND x_counter <= 384 ) OR (x_counter >= 391 AND x_counter <= 400 ) OR (x_counter >= 408 AND x_counter <= 417 ) OR (x_counter >= 441 AND x_counter <= 450 )))
                                        OR ( y_counter = 197 AND ((x_counter >= 177 AND x_counter <= 186 ) OR (x_counter >= 193 AND x_counter <= 202 ) OR (x_counter >= 210 AND x_counter <= 219 ) OR (x_counter >= 226 AND x_counter <= 235 ) OR (x_counter >= 243 AND x_counter <= 252 ) OR (x_counter >= 255 AND x_counter <= 260 ) OR (x_counter >= 263 AND x_counter <= 272 ) OR (x_counter >= 276 AND x_counter <= 285 ) OR (x_counter >= 342 AND x_counter <= 351 ) OR (x_counter >= 358 AND x_counter <= 367 ) OR (x_counter >= 379 AND x_counter <= 396 ) OR (x_counter >= 408 AND x_counter <= 417 ) OR (x_counter >= 441 AND x_counter <= 450 )))
                                        OR ( y_counter = 198 AND ((x_counter >= 177 AND x_counter <= 186 ) OR (x_counter >= 193 AND x_counter <= 202 ) OR (x_counter >= 210 AND x_counter <= 219 ) OR (x_counter >= 226 AND x_counter <= 235 ) OR (x_counter >= 243 AND x_counter <= 252 ) OR (x_counter >= 255 AND x_counter <= 260 ) OR (x_counter >= 263 AND x_counter <= 272 ) OR (x_counter >= 276 AND x_counter <= 285 ) OR (x_counter >= 342 AND x_counter <= 351 ) OR (x_counter >= 358 AND x_counter <= 367 ) OR (x_counter >= 379 AND x_counter <= 396 ) OR (x_counter >= 408 AND x_counter <= 417 ) OR (x_counter >= 441 AND x_counter <= 450 )))
                                        OR ( y_counter = 199 AND ((x_counter >= 177 AND x_counter <= 186 ) OR (x_counter >= 193 AND x_counter <= 202 ) OR (x_counter >= 210 AND x_counter <= 219 ) OR (x_counter >= 226 AND x_counter <= 235 ) OR (x_counter >= 243 AND x_counter <= 252 ) OR (x_counter >= 255 AND x_counter <= 260 ) OR (x_counter >= 263 AND x_counter <= 272 ) OR (x_counter >= 276 AND x_counter <= 285 ) OR (x_counter >= 342 AND x_counter <= 351 ) OR (x_counter >= 358 AND x_counter <= 367 ) OR (x_counter >= 379 AND x_counter <= 396 ) OR (x_counter >= 408 AND x_counter <= 417 ) OR (x_counter >= 441 AND x_counter <= 450 )))
                                        OR ( y_counter = 200 AND ((x_counter >= 177 AND x_counter <= 186 ) OR (x_counter >= 193 AND x_counter <= 202 ) OR (x_counter >= 210 AND x_counter <= 219 ) OR (x_counter >= 226 AND x_counter <= 235 ) OR (x_counter >= 243 AND x_counter <= 252 ) OR (x_counter >= 255 AND x_counter <= 260 ) OR (x_counter >= 263 AND x_counter <= 272 ) OR (x_counter >= 276 AND x_counter <= 285 ) OR (x_counter >= 342 AND x_counter <= 351 ) OR (x_counter >= 358 AND x_counter <= 367 ) OR (x_counter >= 379 AND x_counter <= 396 ) OR (x_counter >= 408 AND x_counter <= 417 ) OR (x_counter >= 441 AND x_counter <= 450 )))
                                        OR ( y_counter = 201 AND ((x_counter >= 181 AND x_counter <= 202 ) OR (x_counter >= 214 AND x_counter <= 235 ) OR (x_counter >= 243 AND x_counter <= 252 ) OR (x_counter >= 263 AND x_counter <= 272 ) OR (x_counter >= 280 AND x_counter <= 297 ) OR (x_counter >= 346 AND x_counter <= 363 ) OR (x_counter >= 383 AND x_counter <= 392 ) OR (x_counter >= 412 AND x_counter <= 429 ) OR (x_counter >= 441 AND x_counter <= 450 )))
                                        OR ( y_counter = 202 AND ((x_counter >= 181 AND x_counter <= 202 ) OR (x_counter >= 214 AND x_counter <= 235 ) OR (x_counter >= 243 AND x_counter <= 252 ) OR (x_counter >= 263 AND x_counter <= 272 ) OR (x_counter >= 280 AND x_counter <= 297 ) OR (x_counter >= 346 AND x_counter <= 363 ) OR (x_counter >= 383 AND x_counter <= 392 ) OR (x_counter >= 412 AND x_counter <= 429 ) OR (x_counter >= 441 AND x_counter <= 450 )))
                                        OR ( y_counter = 203 AND ((x_counter >= 181 AND x_counter <= 202 ) OR (x_counter >= 214 AND x_counter <= 235 ) OR (x_counter >= 243 AND x_counter <= 252 ) OR (x_counter >= 263 AND x_counter <= 272 ) OR (x_counter >= 280 AND x_counter <= 297 ) OR (x_counter >= 346 AND x_counter <= 363 ) OR (x_counter >= 383 AND x_counter <= 392 ) OR (x_counter >= 412 AND x_counter <= 429 ) OR (x_counter >= 441 AND x_counter <= 450 )))
                                        OR ( y_counter = 204 AND ((x_counter >= 181 AND x_counter <= 202 ) OR (x_counter >= 214 AND x_counter <= 235 ) OR (x_counter >= 243 AND x_counter <= 252 ) OR (x_counter >= 263 AND x_counter <= 272 ) OR (x_counter >= 280 AND x_counter <= 297 ) OR (x_counter >= 346 AND x_counter <= 363 ) OR (x_counter >= 383 AND x_counter <= 392 ) OR (x_counter >= 412 AND x_counter <= 429 ) OR (x_counter >= 441 AND x_counter <= 450 )))
                                        OR ( y_counter = 242 AND animation_on ='1' AND ((x_counter >= 409 AND x_counter <= 411 ))) --START ANIMATION
                                        OR ( y_counter = 243 AND animation_on ='1' AND ((x_counter >= 215 AND x_counter <= 220 ) OR (x_counter >= 296 AND x_counter <= 298 ) OR (x_counter >= 312 AND x_counter <= 314 ) OR (x_counter >= 344 AND x_counter <= 346 ) OR (x_counter >= 368 AND x_counter <= 370 ) OR (x_counter >= 409 AND x_counter <= 411 )))
                                        OR ( y_counter = 244 AND animation_on ='1' AND ((x_counter >= 215 AND x_counter <= 217 ) OR (x_counter >= 219 AND x_counter <= 221 ) OR (x_counter >= 296 AND x_counter <= 298 ) OR (x_counter >= 312 AND x_counter <= 314 ) OR (x_counter >= 344 AND x_counter <= 346 ) OR (x_counter >= 368 AND x_counter <= 370 )))
                                        OR ( y_counter = 245 AND animation_on ='1' AND ((x_counter >= 215 AND x_counter <= 217 ) OR (x_counter >= 219 AND x_counter <= 221 ) OR (x_counter >= 223 AND x_counter <= 225 ) OR (x_counter >= 227 AND x_counter <= 229 ) OR (x_counter >= 232 AND x_counter <= 236 ) OR (x_counter >= 240 AND x_counter <= 245 ) OR (x_counter >= 248 AND x_counter <= 253 ) OR (x_counter >= 263 AND x_counter <= 265 ) OR (x_counter >= 267 AND x_counter <= 269 ) OR (x_counter >= 272 AND x_counter <= 276 ) OR (x_counter >= 280 AND x_counter <= 285 ) OR (x_counter >= 288 AND x_counter <= 292 ) OR (x_counter >= 295 AND x_counter <= 301 ) OR (x_counter >= 311 AND x_counter <= 317 ) OR (x_counter >= 320 AND x_counter <= 324 ) OR (x_counter >= 336 AND x_counter <= 341 ) OR (x_counter >= 343 AND x_counter <= 349 ) OR (x_counter >= 352 AND x_counter <= 356 ) OR (x_counter >= 359 AND x_counter <= 361 ) OR (x_counter >= 363 AND x_counter <= 365 ) OR (x_counter >= 367 AND x_counter <= 373 ) OR (x_counter >= 384 AND x_counter <= 388 ) OR (x_counter >= 392 AND x_counter <= 397 ) OR (x_counter >= 400 AND x_counter <= 404 ) OR (x_counter >= 407 AND x_counter <= 411 ) OR (x_counter >= 415 AND x_counter <= 420 )))
                                        OR ( y_counter = 246 AND animation_on ='1' AND ((x_counter >= 215 AND x_counter <= 217 ) OR (x_counter >= 219 AND x_counter <= 221 ) OR (x_counter >= 223 AND x_counter <= 225 ) OR (x_counter >= 226 AND x_counter <= 229 ) OR (x_counter >= 231 AND x_counter <= 233 ) OR (x_counter >= 235 AND x_counter <= 237 ) OR (x_counter >= 239 AND x_counter <= 241 ) OR (x_counter >= 247 AND x_counter <= 249 ) OR (x_counter >= 263 AND x_counter <= 265 ) OR (x_counter >= 266 AND x_counter <= 269 ) OR (x_counter >= 271 AND x_counter <= 273 ) OR (x_counter >= 275 AND x_counter <= 277 ) OR (x_counter >= 279 AND x_counter <= 281 ) OR (x_counter >= 287 AND x_counter <= 289 ) OR (x_counter >= 291 AND x_counter <= 293 ) OR (x_counter >= 296 AND x_counter <= 298 ) OR (x_counter >= 312 AND x_counter <= 314 ) OR (x_counter >= 319 AND x_counter <= 321 ) OR (x_counter >= 323 AND x_counter <= 325 ) OR (x_counter >= 335 AND x_counter <= 337 ) OR (x_counter >= 344 AND x_counter <= 346 ) OR (x_counter >= 355 AND x_counter <= 357 ) OR (x_counter >= 359 AND x_counter <= 361 ) OR (x_counter >= 362 AND x_counter <= 365 ) OR (x_counter >= 368 AND x_counter <= 370 ) OR (x_counter >= 387 AND x_counter <= 389 ) OR (x_counter >= 391 AND x_counter <= 393 ) OR (x_counter >= 395 AND x_counter <= 397 ) OR (x_counter >= 403 AND x_counter <= 405 ) OR (x_counter >= 409 AND x_counter <= 411 ) OR (x_counter >= 415 AND x_counter <= 417 ) OR (x_counter >= 419 AND x_counter <= 421 )))
                                        OR ( y_counter = 247 AND animation_on ='1' AND ((x_counter >= 215 AND x_counter <= 220 ) OR (x_counter >= 223 AND x_counter <= 226 ) OR (x_counter >= 231 AND x_counter <= 233 ) OR (x_counter >= 235 AND x_counter <= 237 ) OR (x_counter >= 239 AND x_counter <= 241 ) OR (x_counter >= 247 AND x_counter <= 249 ) OR (x_counter >= 263 AND x_counter <= 266 ) OR (x_counter >= 271 AND x_counter <= 273 ) OR (x_counter >= 275 AND x_counter <= 277 ) OR (x_counter >= 279 AND x_counter <= 281 ) OR (x_counter >= 287 AND x_counter <= 289 ) OR (x_counter >= 291 AND x_counter <= 293 ) OR (x_counter >= 296 AND x_counter <= 298 ) OR (x_counter >= 312 AND x_counter <= 314 ) OR (x_counter >= 319 AND x_counter <= 321 ) OR (x_counter >= 323 AND x_counter <= 325 ) OR (x_counter >= 335 AND x_counter <= 337 ) OR (x_counter >= 344 AND x_counter <= 346 ) OR (x_counter >= 355 AND x_counter <= 357 ) OR (x_counter >= 359 AND x_counter <= 362 ) OR (x_counter >= 368 AND x_counter <= 370 ) OR (x_counter >= 387 AND x_counter <= 389 ) OR (x_counter >= 391 AND x_counter <= 393 ) OR (x_counter >= 395 AND x_counter <= 397 ) OR (x_counter >= 403 AND x_counter <= 405 ) OR (x_counter >= 409 AND x_counter <= 411 ) OR (x_counter >= 415 AND x_counter <= 417 ) OR (x_counter >= 419 AND x_counter <= 421 )))
                                        OR ( y_counter = 248 AND animation_on ='1' AND ((x_counter >= 215 AND x_counter <= 217 ) OR (x_counter >= 223 AND x_counter <= 225 ) OR (x_counter >= 231 AND x_counter <= 237 ) OR (x_counter >= 240 AND x_counter <= 244 ) OR (x_counter >= 248 AND x_counter <= 252 ) OR (x_counter >= 263 AND x_counter <= 265 ) OR (x_counter >= 271 AND x_counter <= 277 ) OR (x_counter >= 280 AND x_counter <= 284 ) OR (x_counter >= 287 AND x_counter <= 293 ) OR (x_counter >= 296 AND x_counter <= 298 ) OR (x_counter >= 312 AND x_counter <= 314 ) OR (x_counter >= 319 AND x_counter <= 321 ) OR (x_counter >= 323 AND x_counter <= 325 ) OR (x_counter >= 336 AND x_counter <= 340 ) OR (x_counter >= 344 AND x_counter <= 346 ) OR (x_counter >= 352 AND x_counter <= 357 ) OR (x_counter >= 359 AND x_counter <= 361 ) OR (x_counter >= 368 AND x_counter <= 370 ) OR (x_counter >= 384 AND x_counter <= 389 ) OR (x_counter >= 391 AND x_counter <= 393 ) OR (x_counter >= 395 AND x_counter <= 397 ) OR (x_counter >= 400 AND x_counter <= 405 ) OR (x_counter >= 409 AND x_counter <= 411 ) OR (x_counter >= 415 AND x_counter <= 417 ) OR (x_counter >= 419 AND x_counter <= 421 )))
                                        OR ( y_counter = 249 AND animation_on ='1' AND ((x_counter >= 215 AND x_counter <= 217 ) OR (x_counter >= 223 AND x_counter <= 225 ) OR (x_counter >= 231 AND x_counter <= 233 ) OR (x_counter >= 243 AND x_counter <= 245 ) OR (x_counter >= 251 AND x_counter <= 253 ) OR (x_counter >= 263 AND x_counter <= 265 ) OR (x_counter >= 271 AND x_counter <= 273 ) OR (x_counter >= 283 AND x_counter <= 285 ) OR (x_counter >= 287 AND x_counter <= 289 ) OR (x_counter >= 296 AND x_counter <= 298 ) OR (x_counter >= 312 AND x_counter <= 314 ) OR (x_counter >= 319 AND x_counter <= 321 ) OR (x_counter >= 323 AND x_counter <= 325 ) OR (x_counter >= 339 AND x_counter <= 341 ) OR (x_counter >= 344 AND x_counter <= 346 ) OR (x_counter >= 351 AND x_counter <= 353 ) OR (x_counter >= 355 AND x_counter <= 357 ) OR (x_counter >= 359 AND x_counter <= 361 ) OR (x_counter >= 368 AND x_counter <= 370 ) OR (x_counter >= 383 AND x_counter <= 385 ) OR (x_counter >= 387 AND x_counter <= 389 ) OR (x_counter >= 391 AND x_counter <= 393 ) OR (x_counter >= 395 AND x_counter <= 397 ) OR (x_counter >= 399 AND x_counter <= 401 ) OR (x_counter >= 403 AND x_counter <= 405 ) OR (x_counter >= 409 AND x_counter <= 411 ) OR (x_counter >= 415 AND x_counter <= 417 ) OR (x_counter >= 419 AND x_counter <= 421 )))
                                        OR ( y_counter = 250 AND animation_on ='1' AND ((x_counter >= 215 AND x_counter <= 217 ) OR (x_counter >= 223 AND x_counter <= 225 ) OR (x_counter >= 231 AND x_counter <= 233 ) OR (x_counter >= 243 AND x_counter <= 245 ) OR (x_counter >= 251 AND x_counter <= 253 ) OR (x_counter >= 263 AND x_counter <= 265 ) OR (x_counter >= 271 AND x_counter <= 273 ) OR (x_counter >= 283 AND x_counter <= 285 ) OR (x_counter >= 287 AND x_counter <= 289 ) OR (x_counter >= 296 AND x_counter <= 298 ) OR (x_counter >= 312 AND x_counter <= 314 ) OR (x_counter >= 319 AND x_counter <= 321 ) OR (x_counter >= 323 AND x_counter <= 325 ) OR (x_counter >= 339 AND x_counter <= 341 ) OR (x_counter >= 344 AND x_counter <= 346 ) OR (x_counter >= 351 AND x_counter <= 353 ) OR (x_counter >= 355 AND x_counter <= 357 ) OR (x_counter >= 359 AND x_counter <= 361 ) OR (x_counter >= 368 AND x_counter <= 370 ) OR (x_counter >= 383 AND x_counter <= 385 ) OR (x_counter >= 387 AND x_counter <= 389 ) OR (x_counter >= 391 AND x_counter <= 393 ) OR (x_counter >= 395 AND x_counter <= 397 ) OR (x_counter >= 399 AND x_counter <= 401 ) OR (x_counter >= 403 AND x_counter <= 405 ) OR (x_counter >= 409 AND x_counter <= 411 ) OR (x_counter >= 415 AND x_counter <= 417 ) OR (x_counter >= 419 AND x_counter <= 421 )))
                                        OR ( y_counter = 251 AND animation_on ='1' AND ((x_counter >= 215 AND x_counter <= 217 ) OR (x_counter >= 223 AND x_counter <= 225 ) OR (x_counter >= 232 AND x_counter <= 236 ) OR (x_counter >= 239 AND x_counter <= 244 ) OR (x_counter >= 247 AND x_counter <= 252 ) OR (x_counter >= 263 AND x_counter <= 265 ) OR (x_counter >= 272 AND x_counter <= 276 ) OR (x_counter >= 279 AND x_counter <= 284 ) OR (x_counter >= 288 AND x_counter <= 292 ) OR (x_counter >= 297 AND x_counter <= 301 ) OR (x_counter >= 313 AND x_counter <= 317 ) OR (x_counter >= 320 AND x_counter <= 324 ) OR (x_counter >= 335 AND x_counter <= 340 ) OR (x_counter >= 345 AND x_counter <= 349 ) OR (x_counter >= 352 AND x_counter <= 357 ) OR (x_counter >= 359 AND x_counter <= 361 ) OR (x_counter >= 369 AND x_counter <= 373 ) OR (x_counter >= 384 AND x_counter <= 389 ) OR (x_counter >= 392 AND x_counter <= 397 ) OR (x_counter >= 400 AND x_counter <= 405 ) OR (x_counter >= 407 AND x_counter <= 413 ) OR (x_counter >= 415 AND x_counter <= 417 ) OR (x_counter >= 419 AND x_counter <= 421 )))
                                        OR ( y_counter = 252 AND animation_on ='1' AND ((x_counter >= 395 AND x_counter <= 397 )))
                                        OR ( y_counter = 253 AND animation_on ='1' AND ((x_counter >= 395 AND x_counter <= 397 )))
                                        OR ( y_counter = 254 AND animation_on ='1' AND ((x_counter >= 391 AND x_counter <= 396 )))  --END ANIMATION
                                        else "100";

end Behavioral;

